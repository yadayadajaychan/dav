module graphics(
	input vgaclk, // 25 MHz
	input rst, // active low

	input [3:0] grid [0:15],
	input [1:0] state,
	input [9:0] hc,
	input [9:0] vc,

	output reg [11:0] color // RGB
);

	reg bitmap [0:3071];
	reg [11:0] palette [0:23];

	reg [6:0] x;
	reg [6:0] y;
	assign x = hc/7;
	assign y = vc/7;

	reg [3:0] xi;
	reg [3:0] yi;
	assign xi = x % 16;
	assign yi = y % 16;

	reg [3:0] block;
	assign block = x/16 + y/4;

	always @(posedge vgaclk) begin
		if (x >= 64 || y >= 64 || block >= 16) begin
			color <= 12'd0;
		end else begin
			color <= palette[grid[block]*2 + bitmap[grid[block]*256 + xi + yi*16]];
		end
	end

	always @(negedge rst) begin
		bitmap[0] <= 1'b0;
		bitmap[1] <= 1'b0;
		bitmap[2] <= 1'b0;
		bitmap[3] <= 1'b0;
		bitmap[4] <= 1'b0;
		bitmap[5] <= 1'b0;
		bitmap[6] <= 1'b0;
		bitmap[7] <= 1'b0;
		bitmap[8] <= 1'b0;
		bitmap[9] <= 1'b0;
		bitmap[10] <= 1'b0;
		bitmap[11] <= 1'b0;
		bitmap[12] <= 1'b0;
		bitmap[13] <= 1'b0;
		bitmap[14] <= 1'b0;
		bitmap[15] <= 1'b0;
		bitmap[16] <= 1'b0;
		bitmap[17] <= 1'b0;
		bitmap[18] <= 1'b0;
		bitmap[19] <= 1'b0;
		bitmap[20] <= 1'b0;
		bitmap[21] <= 1'b0;
		bitmap[22] <= 1'b0;
		bitmap[23] <= 1'b0;
		bitmap[24] <= 1'b0;
		bitmap[25] <= 1'b0;
		bitmap[26] <= 1'b0;
		bitmap[27] <= 1'b0;
		bitmap[28] <= 1'b0;
		bitmap[29] <= 1'b0;
		bitmap[30] <= 1'b0;
		bitmap[31] <= 1'b0;
		bitmap[32] <= 1'b0;
		bitmap[33] <= 1'b0;
		bitmap[34] <= 1'b0;
		bitmap[35] <= 1'b0;
		bitmap[36] <= 1'b0;
		bitmap[37] <= 1'b0;
		bitmap[38] <= 1'b0;
		bitmap[39] <= 1'b0;
		bitmap[40] <= 1'b0;
		bitmap[41] <= 1'b0;
		bitmap[42] <= 1'b0;
		bitmap[43] <= 1'b0;
		bitmap[44] <= 1'b0;
		bitmap[45] <= 1'b0;
		bitmap[46] <= 1'b0;
		bitmap[47] <= 1'b0;
		bitmap[48] <= 1'b0;
		bitmap[49] <= 1'b0;
		bitmap[50] <= 1'b0;
		bitmap[51] <= 1'b0;
		bitmap[52] <= 1'b0;
		bitmap[53] <= 1'b0;
		bitmap[54] <= 1'b0;
		bitmap[55] <= 1'b0;
		bitmap[56] <= 1'b0;
		bitmap[57] <= 1'b0;
		bitmap[58] <= 1'b0;
		bitmap[59] <= 1'b0;
		bitmap[60] <= 1'b0;
		bitmap[61] <= 1'b0;
		bitmap[62] <= 1'b0;
		bitmap[63] <= 1'b0;
		bitmap[64] <= 1'b0;
		bitmap[65] <= 1'b0;
		bitmap[66] <= 1'b0;
		bitmap[67] <= 1'b0;
		bitmap[68] <= 1'b0;
		bitmap[69] <= 1'b0;
		bitmap[70] <= 1'b0;
		bitmap[71] <= 1'b0;
		bitmap[72] <= 1'b0;
		bitmap[73] <= 1'b0;
		bitmap[74] <= 1'b0;
		bitmap[75] <= 1'b0;
		bitmap[76] <= 1'b0;
		bitmap[77] <= 1'b0;
		bitmap[78] <= 1'b0;
		bitmap[79] <= 1'b0;
		bitmap[80] <= 1'b0;
		bitmap[81] <= 1'b0;
		bitmap[82] <= 1'b0;
		bitmap[83] <= 1'b0;
		bitmap[84] <= 1'b0;
		bitmap[85] <= 1'b0;
		bitmap[86] <= 1'b0;
		bitmap[87] <= 1'b0;
		bitmap[88] <= 1'b0;
		bitmap[89] <= 1'b0;
		bitmap[90] <= 1'b0;
		bitmap[91] <= 1'b0;
		bitmap[92] <= 1'b0;
		bitmap[93] <= 1'b0;
		bitmap[94] <= 1'b0;
		bitmap[95] <= 1'b0;
		bitmap[96] <= 1'b0;
		bitmap[97] <= 1'b0;
		bitmap[98] <= 1'b0;
		bitmap[99] <= 1'b0;
		bitmap[100] <= 1'b0;
		bitmap[101] <= 1'b0;
		bitmap[102] <= 1'b0;
		bitmap[103] <= 1'b0;
		bitmap[104] <= 1'b0;
		bitmap[105] <= 1'b0;
		bitmap[106] <= 1'b0;
		bitmap[107] <= 1'b0;
		bitmap[108] <= 1'b0;
		bitmap[109] <= 1'b0;
		bitmap[110] <= 1'b0;
		bitmap[111] <= 1'b0;
		bitmap[112] <= 1'b0;
		bitmap[113] <= 1'b0;
		bitmap[114] <= 1'b0;
		bitmap[115] <= 1'b0;
		bitmap[116] <= 1'b0;
		bitmap[117] <= 1'b0;
		bitmap[118] <= 1'b0;
		bitmap[119] <= 1'b0;
		bitmap[120] <= 1'b0;
		bitmap[121] <= 1'b0;
		bitmap[122] <= 1'b0;
		bitmap[123] <= 1'b0;
		bitmap[124] <= 1'b0;
		bitmap[125] <= 1'b0;
		bitmap[126] <= 1'b0;
		bitmap[127] <= 1'b0;
		bitmap[128] <= 1'b0;
		bitmap[129] <= 1'b0;
		bitmap[130] <= 1'b0;
		bitmap[131] <= 1'b0;
		bitmap[132] <= 1'b0;
		bitmap[133] <= 1'b0;
		bitmap[134] <= 1'b0;
		bitmap[135] <= 1'b0;
		bitmap[136] <= 1'b0;
		bitmap[137] <= 1'b0;
		bitmap[138] <= 1'b0;
		bitmap[139] <= 1'b0;
		bitmap[140] <= 1'b0;
		bitmap[141] <= 1'b0;
		bitmap[142] <= 1'b0;
		bitmap[143] <= 1'b0;
		bitmap[144] <= 1'b0;
		bitmap[145] <= 1'b0;
		bitmap[146] <= 1'b0;
		bitmap[147] <= 1'b0;
		bitmap[148] <= 1'b0;
		bitmap[149] <= 1'b0;
		bitmap[150] <= 1'b0;
		bitmap[151] <= 1'b0;
		bitmap[152] <= 1'b0;
		bitmap[153] <= 1'b0;
		bitmap[154] <= 1'b0;
		bitmap[155] <= 1'b0;
		bitmap[156] <= 1'b0;
		bitmap[157] <= 1'b0;
		bitmap[158] <= 1'b0;
		bitmap[159] <= 1'b0;
		bitmap[160] <= 1'b0;
		bitmap[161] <= 1'b0;
		bitmap[162] <= 1'b0;
		bitmap[163] <= 1'b0;
		bitmap[164] <= 1'b0;
		bitmap[165] <= 1'b0;
		bitmap[166] <= 1'b0;
		bitmap[167] <= 1'b0;
		bitmap[168] <= 1'b0;
		bitmap[169] <= 1'b0;
		bitmap[170] <= 1'b0;
		bitmap[171] <= 1'b0;
		bitmap[172] <= 1'b0;
		bitmap[173] <= 1'b0;
		bitmap[174] <= 1'b0;
		bitmap[175] <= 1'b0;
		bitmap[176] <= 1'b0;
		bitmap[177] <= 1'b0;
		bitmap[178] <= 1'b0;
		bitmap[179] <= 1'b0;
		bitmap[180] <= 1'b0;
		bitmap[181] <= 1'b0;
		bitmap[182] <= 1'b0;
		bitmap[183] <= 1'b0;
		bitmap[184] <= 1'b0;
		bitmap[185] <= 1'b0;
		bitmap[186] <= 1'b0;
		bitmap[187] <= 1'b0;
		bitmap[188] <= 1'b0;
		bitmap[189] <= 1'b0;
		bitmap[190] <= 1'b0;
		bitmap[191] <= 1'b0;
		bitmap[192] <= 1'b0;
		bitmap[193] <= 1'b0;
		bitmap[194] <= 1'b0;
		bitmap[195] <= 1'b0;
		bitmap[196] <= 1'b0;
		bitmap[197] <= 1'b0;
		bitmap[198] <= 1'b0;
		bitmap[199] <= 1'b0;
		bitmap[200] <= 1'b0;
		bitmap[201] <= 1'b0;
		bitmap[202] <= 1'b0;
		bitmap[203] <= 1'b0;
		bitmap[204] <= 1'b0;
		bitmap[205] <= 1'b0;
		bitmap[206] <= 1'b0;
		bitmap[207] <= 1'b0;
		bitmap[208] <= 1'b0;
		bitmap[209] <= 1'b0;
		bitmap[210] <= 1'b0;
		bitmap[211] <= 1'b0;
		bitmap[212] <= 1'b0;
		bitmap[213] <= 1'b0;
		bitmap[214] <= 1'b0;
		bitmap[215] <= 1'b0;
		bitmap[216] <= 1'b0;
		bitmap[217] <= 1'b0;
		bitmap[218] <= 1'b0;
		bitmap[219] <= 1'b0;
		bitmap[220] <= 1'b0;
		bitmap[221] <= 1'b0;
		bitmap[222] <= 1'b0;
		bitmap[223] <= 1'b0;
		bitmap[224] <= 1'b0;
		bitmap[225] <= 1'b0;
		bitmap[226] <= 1'b0;
		bitmap[227] <= 1'b0;
		bitmap[228] <= 1'b0;
		bitmap[229] <= 1'b0;
		bitmap[230] <= 1'b0;
		bitmap[231] <= 1'b0;
		bitmap[232] <= 1'b0;
		bitmap[233] <= 1'b0;
		bitmap[234] <= 1'b0;
		bitmap[235] <= 1'b0;
		bitmap[236] <= 1'b0;
		bitmap[237] <= 1'b0;
		bitmap[238] <= 1'b0;
		bitmap[239] <= 1'b0;
		bitmap[240] <= 1'b0;
		bitmap[241] <= 1'b0;
		bitmap[242] <= 1'b0;
		bitmap[243] <= 1'b0;
		bitmap[244] <= 1'b0;
		bitmap[245] <= 1'b0;
		bitmap[246] <= 1'b0;
		bitmap[247] <= 1'b0;
		bitmap[248] <= 1'b0;
		bitmap[249] <= 1'b0;
		bitmap[250] <= 1'b0;
		bitmap[251] <= 1'b0;
		bitmap[252] <= 1'b0;
		bitmap[253] <= 1'b0;
		bitmap[254] <= 1'b0;
		bitmap[255] <= 1'b0;
		bitmap[256] <= 1'b0;
		bitmap[257] <= 1'b0;
		bitmap[258] <= 1'b0;
		bitmap[259] <= 1'b0;
		bitmap[260] <= 1'b0;
		bitmap[261] <= 1'b0;
		bitmap[262] <= 1'b0;
		bitmap[263] <= 1'b0;
		bitmap[264] <= 1'b0;
		bitmap[265] <= 1'b0;
		bitmap[266] <= 1'b0;
		bitmap[267] <= 1'b0;
		bitmap[268] <= 1'b0;
		bitmap[269] <= 1'b0;
		bitmap[270] <= 1'b0;
		bitmap[271] <= 1'b0;
		bitmap[272] <= 1'b0;
		bitmap[273] <= 1'b0;
		bitmap[274] <= 1'b0;
		bitmap[275] <= 1'b1;
		bitmap[276] <= 1'b1;
		bitmap[277] <= 1'b0;
		bitmap[278] <= 1'b0;
		bitmap[279] <= 1'b0;
		bitmap[280] <= 1'b0;
		bitmap[281] <= 1'b0;
		bitmap[282] <= 1'b0;
		bitmap[283] <= 1'b0;
		bitmap[284] <= 1'b0;
		bitmap[285] <= 1'b0;
		bitmap[286] <= 1'b0;
		bitmap[287] <= 1'b0;
		bitmap[288] <= 1'b0;
		bitmap[289] <= 1'b0;
		bitmap[290] <= 1'b1;
		bitmap[291] <= 1'b0;
		bitmap[292] <= 1'b0;
		bitmap[293] <= 1'b1;
		bitmap[294] <= 1'b0;
		bitmap[295] <= 1'b0;
		bitmap[296] <= 1'b0;
		bitmap[297] <= 1'b0;
		bitmap[298] <= 1'b0;
		bitmap[299] <= 1'b0;
		bitmap[300] <= 1'b0;
		bitmap[301] <= 1'b0;
		bitmap[302] <= 1'b0;
		bitmap[303] <= 1'b0;
		bitmap[304] <= 1'b0;
		bitmap[305] <= 1'b0;
		bitmap[306] <= 1'b0;
		bitmap[307] <= 1'b0;
		bitmap[308] <= 1'b0;
		bitmap[309] <= 1'b1;
		bitmap[310] <= 1'b0;
		bitmap[311] <= 1'b0;
		bitmap[312] <= 1'b0;
		bitmap[313] <= 1'b0;
		bitmap[314] <= 1'b0;
		bitmap[315] <= 1'b0;
		bitmap[316] <= 1'b0;
		bitmap[317] <= 1'b0;
		bitmap[318] <= 1'b0;
		bitmap[319] <= 1'b0;
		bitmap[320] <= 1'b0;
		bitmap[321] <= 1'b0;
		bitmap[322] <= 1'b0;
		bitmap[323] <= 1'b0;
		bitmap[324] <= 1'b1;
		bitmap[325] <= 1'b0;
		bitmap[326] <= 1'b0;
		bitmap[327] <= 1'b0;
		bitmap[328] <= 1'b0;
		bitmap[329] <= 1'b0;
		bitmap[330] <= 1'b0;
		bitmap[331] <= 1'b0;
		bitmap[332] <= 1'b0;
		bitmap[333] <= 1'b0;
		bitmap[334] <= 1'b0;
		bitmap[335] <= 1'b0;
		bitmap[336] <= 1'b0;
		bitmap[337] <= 1'b0;
		bitmap[338] <= 1'b0;
		bitmap[339] <= 1'b1;
		bitmap[340] <= 1'b0;
		bitmap[341] <= 1'b0;
		bitmap[342] <= 1'b0;
		bitmap[343] <= 1'b0;
		bitmap[344] <= 1'b0;
		bitmap[345] <= 1'b0;
		bitmap[346] <= 1'b0;
		bitmap[347] <= 1'b0;
		bitmap[348] <= 1'b0;
		bitmap[349] <= 1'b0;
		bitmap[350] <= 1'b0;
		bitmap[351] <= 1'b0;
		bitmap[352] <= 1'b0;
		bitmap[353] <= 1'b0;
		bitmap[354] <= 1'b1;
		bitmap[355] <= 1'b1;
		bitmap[356] <= 1'b1;
		bitmap[357] <= 1'b1;
		bitmap[358] <= 1'b0;
		bitmap[359] <= 1'b0;
		bitmap[360] <= 1'b0;
		bitmap[361] <= 1'b0;
		bitmap[362] <= 1'b0;
		bitmap[363] <= 1'b0;
		bitmap[364] <= 1'b0;
		bitmap[365] <= 1'b0;
		bitmap[366] <= 1'b0;
		bitmap[367] <= 1'b0;
		bitmap[368] <= 1'b0;
		bitmap[369] <= 1'b0;
		bitmap[370] <= 1'b0;
		bitmap[371] <= 1'b0;
		bitmap[372] <= 1'b0;
		bitmap[373] <= 1'b0;
		bitmap[374] <= 1'b0;
		bitmap[375] <= 1'b0;
		bitmap[376] <= 1'b0;
		bitmap[377] <= 1'b0;
		bitmap[378] <= 1'b0;
		bitmap[379] <= 1'b0;
		bitmap[380] <= 1'b0;
		bitmap[381] <= 1'b0;
		bitmap[382] <= 1'b0;
		bitmap[383] <= 1'b0;
		bitmap[384] <= 1'b0;
		bitmap[385] <= 1'b0;
		bitmap[386] <= 1'b0;
		bitmap[387] <= 1'b0;
		bitmap[388] <= 1'b0;
		bitmap[389] <= 1'b0;
		bitmap[390] <= 1'b0;
		bitmap[391] <= 1'b0;
		bitmap[392] <= 1'b0;
		bitmap[393] <= 1'b0;
		bitmap[394] <= 1'b0;
		bitmap[395] <= 1'b0;
		bitmap[396] <= 1'b0;
		bitmap[397] <= 1'b0;
		bitmap[398] <= 1'b0;
		bitmap[399] <= 1'b0;
		bitmap[400] <= 1'b0;
		bitmap[401] <= 1'b0;
		bitmap[402] <= 1'b0;
		bitmap[403] <= 1'b0;
		bitmap[404] <= 1'b0;
		bitmap[405] <= 1'b0;
		bitmap[406] <= 1'b0;
		bitmap[407] <= 1'b0;
		bitmap[408] <= 1'b0;
		bitmap[409] <= 1'b0;
		bitmap[410] <= 1'b0;
		bitmap[411] <= 1'b0;
		bitmap[412] <= 1'b0;
		bitmap[413] <= 1'b0;
		bitmap[414] <= 1'b0;
		bitmap[415] <= 1'b0;
		bitmap[416] <= 1'b0;
		bitmap[417] <= 1'b0;
		bitmap[418] <= 1'b0;
		bitmap[419] <= 1'b0;
		bitmap[420] <= 1'b0;
		bitmap[421] <= 1'b0;
		bitmap[422] <= 1'b0;
		bitmap[423] <= 1'b0;
		bitmap[424] <= 1'b0;
		bitmap[425] <= 1'b0;
		bitmap[426] <= 1'b0;
		bitmap[427] <= 1'b0;
		bitmap[428] <= 1'b0;
		bitmap[429] <= 1'b0;
		bitmap[430] <= 1'b0;
		bitmap[431] <= 1'b0;
		bitmap[432] <= 1'b0;
		bitmap[433] <= 1'b0;
		bitmap[434] <= 1'b0;
		bitmap[435] <= 1'b0;
		bitmap[436] <= 1'b0;
		bitmap[437] <= 1'b0;
		bitmap[438] <= 1'b0;
		bitmap[439] <= 1'b0;
		bitmap[440] <= 1'b0;
		bitmap[441] <= 1'b0;
		bitmap[442] <= 1'b0;
		bitmap[443] <= 1'b0;
		bitmap[444] <= 1'b0;
		bitmap[445] <= 1'b0;
		bitmap[446] <= 1'b0;
		bitmap[447] <= 1'b0;
		bitmap[448] <= 1'b0;
		bitmap[449] <= 1'b0;
		bitmap[450] <= 1'b0;
		bitmap[451] <= 1'b0;
		bitmap[452] <= 1'b0;
		bitmap[453] <= 1'b0;
		bitmap[454] <= 1'b0;
		bitmap[455] <= 1'b0;
		bitmap[456] <= 1'b0;
		bitmap[457] <= 1'b0;
		bitmap[458] <= 1'b0;
		bitmap[459] <= 1'b0;
		bitmap[460] <= 1'b0;
		bitmap[461] <= 1'b0;
		bitmap[462] <= 1'b0;
		bitmap[463] <= 1'b0;
		bitmap[464] <= 1'b0;
		bitmap[465] <= 1'b0;
		bitmap[466] <= 1'b0;
		bitmap[467] <= 1'b0;
		bitmap[468] <= 1'b0;
		bitmap[469] <= 1'b0;
		bitmap[470] <= 1'b0;
		bitmap[471] <= 1'b0;
		bitmap[472] <= 1'b0;
		bitmap[473] <= 1'b0;
		bitmap[474] <= 1'b0;
		bitmap[475] <= 1'b0;
		bitmap[476] <= 1'b0;
		bitmap[477] <= 1'b0;
		bitmap[478] <= 1'b0;
		bitmap[479] <= 1'b0;
		bitmap[480] <= 1'b0;
		bitmap[481] <= 1'b0;
		bitmap[482] <= 1'b0;
		bitmap[483] <= 1'b0;
		bitmap[484] <= 1'b0;
		bitmap[485] <= 1'b0;
		bitmap[486] <= 1'b0;
		bitmap[487] <= 1'b0;
		bitmap[488] <= 1'b0;
		bitmap[489] <= 1'b0;
		bitmap[490] <= 1'b0;
		bitmap[491] <= 1'b0;
		bitmap[492] <= 1'b0;
		bitmap[493] <= 1'b0;
		bitmap[494] <= 1'b0;
		bitmap[495] <= 1'b0;
		bitmap[496] <= 1'b0;
		bitmap[497] <= 1'b0;
		bitmap[498] <= 1'b0;
		bitmap[499] <= 1'b0;
		bitmap[500] <= 1'b0;
		bitmap[501] <= 1'b0;
		bitmap[502] <= 1'b0;
		bitmap[503] <= 1'b0;
		bitmap[504] <= 1'b0;
		bitmap[505] <= 1'b0;
		bitmap[506] <= 1'b0;
		bitmap[507] <= 1'b0;
		bitmap[508] <= 1'b0;
		bitmap[509] <= 1'b0;
		bitmap[510] <= 1'b0;
		bitmap[511] <= 1'b0;
		bitmap[512] <= 1'b0;
		bitmap[513] <= 1'b0;
		bitmap[514] <= 1'b0;
		bitmap[515] <= 1'b0;
		bitmap[516] <= 1'b0;
		bitmap[517] <= 1'b0;
		bitmap[518] <= 1'b0;
		bitmap[519] <= 1'b0;
		bitmap[520] <= 1'b0;
		bitmap[521] <= 1'b0;
		bitmap[522] <= 1'b0;
		bitmap[523] <= 1'b0;
		bitmap[524] <= 1'b0;
		bitmap[525] <= 1'b0;
		bitmap[526] <= 1'b0;
		bitmap[527] <= 1'b0;
		bitmap[528] <= 1'b0;
		bitmap[529] <= 1'b0;
		bitmap[530] <= 1'b0;
		bitmap[531] <= 1'b0;
		bitmap[532] <= 1'b1;
		bitmap[533] <= 1'b1;
		bitmap[534] <= 1'b0;
		bitmap[535] <= 1'b0;
		bitmap[536] <= 1'b0;
		bitmap[537] <= 1'b0;
		bitmap[538] <= 1'b0;
		bitmap[539] <= 1'b0;
		bitmap[540] <= 1'b0;
		bitmap[541] <= 1'b0;
		bitmap[542] <= 1'b0;
		bitmap[543] <= 1'b0;
		bitmap[544] <= 1'b0;
		bitmap[545] <= 1'b0;
		bitmap[546] <= 1'b0;
		bitmap[547] <= 1'b1;
		bitmap[548] <= 1'b0;
		bitmap[549] <= 1'b1;
		bitmap[550] <= 1'b0;
		bitmap[551] <= 1'b0;
		bitmap[552] <= 1'b0;
		bitmap[553] <= 1'b0;
		bitmap[554] <= 1'b0;
		bitmap[555] <= 1'b0;
		bitmap[556] <= 1'b0;
		bitmap[557] <= 1'b0;
		bitmap[558] <= 1'b0;
		bitmap[559] <= 1'b0;
		bitmap[560] <= 1'b0;
		bitmap[561] <= 1'b0;
		bitmap[562] <= 1'b1;
		bitmap[563] <= 1'b0;
		bitmap[564] <= 1'b0;
		bitmap[565] <= 1'b1;
		bitmap[566] <= 1'b0;
		bitmap[567] <= 1'b0;
		bitmap[568] <= 1'b0;
		bitmap[569] <= 1'b0;
		bitmap[570] <= 1'b0;
		bitmap[571] <= 1'b0;
		bitmap[572] <= 1'b0;
		bitmap[573] <= 1'b0;
		bitmap[574] <= 1'b0;
		bitmap[575] <= 1'b0;
		bitmap[576] <= 1'b0;
		bitmap[577] <= 1'b0;
		bitmap[578] <= 1'b1;
		bitmap[579] <= 1'b1;
		bitmap[580] <= 1'b1;
		bitmap[581] <= 1'b1;
		bitmap[582] <= 1'b1;
		bitmap[583] <= 1'b0;
		bitmap[584] <= 1'b0;
		bitmap[585] <= 1'b0;
		bitmap[586] <= 1'b0;
		bitmap[587] <= 1'b0;
		bitmap[588] <= 1'b0;
		bitmap[589] <= 1'b0;
		bitmap[590] <= 1'b0;
		bitmap[591] <= 1'b0;
		bitmap[592] <= 1'b0;
		bitmap[593] <= 1'b0;
		bitmap[594] <= 1'b0;
		bitmap[595] <= 1'b0;
		bitmap[596] <= 1'b0;
		bitmap[597] <= 1'b1;
		bitmap[598] <= 1'b0;
		bitmap[599] <= 1'b0;
		bitmap[600] <= 1'b0;
		bitmap[601] <= 1'b0;
		bitmap[602] <= 1'b0;
		bitmap[603] <= 1'b0;
		bitmap[604] <= 1'b0;
		bitmap[605] <= 1'b0;
		bitmap[606] <= 1'b0;
		bitmap[607] <= 1'b0;
		bitmap[608] <= 1'b0;
		bitmap[609] <= 1'b0;
		bitmap[610] <= 1'b0;
		bitmap[611] <= 1'b0;
		bitmap[612] <= 1'b0;
		bitmap[613] <= 1'b1;
		bitmap[614] <= 1'b0;
		bitmap[615] <= 1'b0;
		bitmap[616] <= 1'b0;
		bitmap[617] <= 1'b0;
		bitmap[618] <= 1'b0;
		bitmap[619] <= 1'b0;
		bitmap[620] <= 1'b0;
		bitmap[621] <= 1'b0;
		bitmap[622] <= 1'b0;
		bitmap[623] <= 1'b0;
		bitmap[624] <= 1'b0;
		bitmap[625] <= 1'b0;
		bitmap[626] <= 1'b0;
		bitmap[627] <= 1'b0;
		bitmap[628] <= 1'b0;
		bitmap[629] <= 1'b0;
		bitmap[630] <= 1'b0;
		bitmap[631] <= 1'b0;
		bitmap[632] <= 1'b0;
		bitmap[633] <= 1'b0;
		bitmap[634] <= 1'b0;
		bitmap[635] <= 1'b0;
		bitmap[636] <= 1'b0;
		bitmap[637] <= 1'b0;
		bitmap[638] <= 1'b0;
		bitmap[639] <= 1'b0;
		bitmap[640] <= 1'b0;
		bitmap[641] <= 1'b0;
		bitmap[642] <= 1'b0;
		bitmap[643] <= 1'b0;
		bitmap[644] <= 1'b0;
		bitmap[645] <= 1'b0;
		bitmap[646] <= 1'b0;
		bitmap[647] <= 1'b0;
		bitmap[648] <= 1'b0;
		bitmap[649] <= 1'b0;
		bitmap[650] <= 1'b0;
		bitmap[651] <= 1'b0;
		bitmap[652] <= 1'b0;
		bitmap[653] <= 1'b0;
		bitmap[654] <= 1'b0;
		bitmap[655] <= 1'b0;
		bitmap[656] <= 1'b0;
		bitmap[657] <= 1'b0;
		bitmap[658] <= 1'b0;
		bitmap[659] <= 1'b0;
		bitmap[660] <= 1'b0;
		bitmap[661] <= 1'b0;
		bitmap[662] <= 1'b0;
		bitmap[663] <= 1'b0;
		bitmap[664] <= 1'b0;
		bitmap[665] <= 1'b0;
		bitmap[666] <= 1'b0;
		bitmap[667] <= 1'b0;
		bitmap[668] <= 1'b0;
		bitmap[669] <= 1'b0;
		bitmap[670] <= 1'b0;
		bitmap[671] <= 1'b0;
		bitmap[672] <= 1'b0;
		bitmap[673] <= 1'b0;
		bitmap[674] <= 1'b0;
		bitmap[675] <= 1'b0;
		bitmap[676] <= 1'b0;
		bitmap[677] <= 1'b0;
		bitmap[678] <= 1'b0;
		bitmap[679] <= 1'b0;
		bitmap[680] <= 1'b0;
		bitmap[681] <= 1'b0;
		bitmap[682] <= 1'b0;
		bitmap[683] <= 1'b0;
		bitmap[684] <= 1'b0;
		bitmap[685] <= 1'b0;
		bitmap[686] <= 1'b0;
		bitmap[687] <= 1'b0;
		bitmap[688] <= 1'b0;
		bitmap[689] <= 1'b0;
		bitmap[690] <= 1'b0;
		bitmap[691] <= 1'b0;
		bitmap[692] <= 1'b0;
		bitmap[693] <= 1'b0;
		bitmap[694] <= 1'b0;
		bitmap[695] <= 1'b0;
		bitmap[696] <= 1'b0;
		bitmap[697] <= 1'b0;
		bitmap[698] <= 1'b0;
		bitmap[699] <= 1'b0;
		bitmap[700] <= 1'b0;
		bitmap[701] <= 1'b0;
		bitmap[702] <= 1'b0;
		bitmap[703] <= 1'b0;
		bitmap[704] <= 1'b0;
		bitmap[705] <= 1'b0;
		bitmap[706] <= 1'b0;
		bitmap[707] <= 1'b0;
		bitmap[708] <= 1'b0;
		bitmap[709] <= 1'b0;
		bitmap[710] <= 1'b0;
		bitmap[711] <= 1'b0;
		bitmap[712] <= 1'b0;
		bitmap[713] <= 1'b0;
		bitmap[714] <= 1'b0;
		bitmap[715] <= 1'b0;
		bitmap[716] <= 1'b0;
		bitmap[717] <= 1'b0;
		bitmap[718] <= 1'b0;
		bitmap[719] <= 1'b0;
		bitmap[720] <= 1'b0;
		bitmap[721] <= 1'b0;
		bitmap[722] <= 1'b0;
		bitmap[723] <= 1'b0;
		bitmap[724] <= 1'b0;
		bitmap[725] <= 1'b0;
		bitmap[726] <= 1'b0;
		bitmap[727] <= 1'b0;
		bitmap[728] <= 1'b0;
		bitmap[729] <= 1'b0;
		bitmap[730] <= 1'b0;
		bitmap[731] <= 1'b0;
		bitmap[732] <= 1'b0;
		bitmap[733] <= 1'b0;
		bitmap[734] <= 1'b0;
		bitmap[735] <= 1'b0;
		bitmap[736] <= 1'b0;
		bitmap[737] <= 1'b0;
		bitmap[738] <= 1'b0;
		bitmap[739] <= 1'b0;
		bitmap[740] <= 1'b0;
		bitmap[741] <= 1'b0;
		bitmap[742] <= 1'b0;
		bitmap[743] <= 1'b0;
		bitmap[744] <= 1'b0;
		bitmap[745] <= 1'b0;
		bitmap[746] <= 1'b0;
		bitmap[747] <= 1'b0;
		bitmap[748] <= 1'b0;
		bitmap[749] <= 1'b0;
		bitmap[750] <= 1'b0;
		bitmap[751] <= 1'b0;
		bitmap[752] <= 1'b0;
		bitmap[753] <= 1'b0;
		bitmap[754] <= 1'b0;
		bitmap[755] <= 1'b0;
		bitmap[756] <= 1'b0;
		bitmap[757] <= 1'b0;
		bitmap[758] <= 1'b0;
		bitmap[759] <= 1'b0;
		bitmap[760] <= 1'b0;
		bitmap[761] <= 1'b0;
		bitmap[762] <= 1'b0;
		bitmap[763] <= 1'b0;
		bitmap[764] <= 1'b0;
		bitmap[765] <= 1'b0;
		bitmap[766] <= 1'b0;
		bitmap[767] <= 1'b0;
		bitmap[768] <= 1'b0;
		bitmap[769] <= 1'b0;
		bitmap[770] <= 1'b0;
		bitmap[771] <= 1'b0;
		bitmap[772] <= 1'b0;
		bitmap[773] <= 1'b0;
		bitmap[774] <= 1'b0;
		bitmap[775] <= 1'b0;
		bitmap[776] <= 1'b0;
		bitmap[777] <= 1'b0;
		bitmap[778] <= 1'b0;
		bitmap[779] <= 1'b0;
		bitmap[780] <= 1'b0;
		bitmap[781] <= 1'b0;
		bitmap[782] <= 1'b0;
		bitmap[783] <= 1'b0;
		bitmap[784] <= 1'b0;
		bitmap[785] <= 1'b0;
		bitmap[786] <= 1'b1;
		bitmap[787] <= 1'b1;
		bitmap[788] <= 1'b1;
		bitmap[789] <= 1'b1;
		bitmap[790] <= 1'b0;
		bitmap[791] <= 1'b0;
		bitmap[792] <= 1'b0;
		bitmap[793] <= 1'b0;
		bitmap[794] <= 1'b0;
		bitmap[795] <= 1'b0;
		bitmap[796] <= 1'b0;
		bitmap[797] <= 1'b0;
		bitmap[798] <= 1'b0;
		bitmap[799] <= 1'b0;
		bitmap[800] <= 1'b0;
		bitmap[801] <= 1'b0;
		bitmap[802] <= 1'b1;
		bitmap[803] <= 1'b0;
		bitmap[804] <= 1'b0;
		bitmap[805] <= 1'b1;
		bitmap[806] <= 1'b0;
		bitmap[807] <= 1'b0;
		bitmap[808] <= 1'b0;
		bitmap[809] <= 1'b0;
		bitmap[810] <= 1'b0;
		bitmap[811] <= 1'b0;
		bitmap[812] <= 1'b0;
		bitmap[813] <= 1'b0;
		bitmap[814] <= 1'b0;
		bitmap[815] <= 1'b0;
		bitmap[816] <= 1'b0;
		bitmap[817] <= 1'b0;
		bitmap[818] <= 1'b1;
		bitmap[819] <= 1'b0;
		bitmap[820] <= 1'b0;
		bitmap[821] <= 1'b1;
		bitmap[822] <= 1'b0;
		bitmap[823] <= 1'b0;
		bitmap[824] <= 1'b0;
		bitmap[825] <= 1'b0;
		bitmap[826] <= 1'b0;
		bitmap[827] <= 1'b0;
		bitmap[828] <= 1'b0;
		bitmap[829] <= 1'b0;
		bitmap[830] <= 1'b0;
		bitmap[831] <= 1'b0;
		bitmap[832] <= 1'b0;
		bitmap[833] <= 1'b0;
		bitmap[834] <= 1'b1;
		bitmap[835] <= 1'b1;
		bitmap[836] <= 1'b1;
		bitmap[837] <= 1'b1;
		bitmap[838] <= 1'b0;
		bitmap[839] <= 1'b0;
		bitmap[840] <= 1'b0;
		bitmap[841] <= 1'b0;
		bitmap[842] <= 1'b0;
		bitmap[843] <= 1'b0;
		bitmap[844] <= 1'b0;
		bitmap[845] <= 1'b0;
		bitmap[846] <= 1'b0;
		bitmap[847] <= 1'b0;
		bitmap[848] <= 1'b0;
		bitmap[849] <= 1'b0;
		bitmap[850] <= 1'b1;
		bitmap[851] <= 1'b0;
		bitmap[852] <= 1'b0;
		bitmap[853] <= 1'b1;
		bitmap[854] <= 1'b0;
		bitmap[855] <= 1'b0;
		bitmap[856] <= 1'b0;
		bitmap[857] <= 1'b0;
		bitmap[858] <= 1'b0;
		bitmap[859] <= 1'b0;
		bitmap[860] <= 1'b0;
		bitmap[861] <= 1'b0;
		bitmap[862] <= 1'b0;
		bitmap[863] <= 1'b0;
		bitmap[864] <= 1'b0;
		bitmap[865] <= 1'b0;
		bitmap[866] <= 1'b1;
		bitmap[867] <= 1'b1;
		bitmap[868] <= 1'b1;
		bitmap[869] <= 1'b1;
		bitmap[870] <= 1'b0;
		bitmap[871] <= 1'b0;
		bitmap[872] <= 1'b0;
		bitmap[873] <= 1'b0;
		bitmap[874] <= 1'b0;
		bitmap[875] <= 1'b0;
		bitmap[876] <= 1'b0;
		bitmap[877] <= 1'b0;
		bitmap[878] <= 1'b0;
		bitmap[879] <= 1'b0;
		bitmap[880] <= 1'b0;
		bitmap[881] <= 1'b0;
		bitmap[882] <= 1'b0;
		bitmap[883] <= 1'b0;
		bitmap[884] <= 1'b0;
		bitmap[885] <= 1'b0;
		bitmap[886] <= 1'b0;
		bitmap[887] <= 1'b0;
		bitmap[888] <= 1'b0;
		bitmap[889] <= 1'b0;
		bitmap[890] <= 1'b0;
		bitmap[891] <= 1'b0;
		bitmap[892] <= 1'b0;
		bitmap[893] <= 1'b0;
		bitmap[894] <= 1'b0;
		bitmap[895] <= 1'b0;
		bitmap[896] <= 1'b0;
		bitmap[897] <= 1'b0;
		bitmap[898] <= 1'b0;
		bitmap[899] <= 1'b0;
		bitmap[900] <= 1'b0;
		bitmap[901] <= 1'b0;
		bitmap[902] <= 1'b0;
		bitmap[903] <= 1'b0;
		bitmap[904] <= 1'b0;
		bitmap[905] <= 1'b0;
		bitmap[906] <= 1'b0;
		bitmap[907] <= 1'b0;
		bitmap[908] <= 1'b0;
		bitmap[909] <= 1'b0;
		bitmap[910] <= 1'b0;
		bitmap[911] <= 1'b0;
		bitmap[912] <= 1'b0;
		bitmap[913] <= 1'b0;
		bitmap[914] <= 1'b0;
		bitmap[915] <= 1'b0;
		bitmap[916] <= 1'b0;
		bitmap[917] <= 1'b0;
		bitmap[918] <= 1'b0;
		bitmap[919] <= 1'b0;
		bitmap[920] <= 1'b0;
		bitmap[921] <= 1'b0;
		bitmap[922] <= 1'b0;
		bitmap[923] <= 1'b0;
		bitmap[924] <= 1'b0;
		bitmap[925] <= 1'b0;
		bitmap[926] <= 1'b0;
		bitmap[927] <= 1'b0;
		bitmap[928] <= 1'b0;
		bitmap[929] <= 1'b0;
		bitmap[930] <= 1'b0;
		bitmap[931] <= 1'b0;
		bitmap[932] <= 1'b0;
		bitmap[933] <= 1'b0;
		bitmap[934] <= 1'b0;
		bitmap[935] <= 1'b0;
		bitmap[936] <= 1'b0;
		bitmap[937] <= 1'b0;
		bitmap[938] <= 1'b0;
		bitmap[939] <= 1'b0;
		bitmap[940] <= 1'b0;
		bitmap[941] <= 1'b0;
		bitmap[942] <= 1'b0;
		bitmap[943] <= 1'b0;
		bitmap[944] <= 1'b0;
		bitmap[945] <= 1'b0;
		bitmap[946] <= 1'b0;
		bitmap[947] <= 1'b0;
		bitmap[948] <= 1'b0;
		bitmap[949] <= 1'b0;
		bitmap[950] <= 1'b0;
		bitmap[951] <= 1'b0;
		bitmap[952] <= 1'b0;
		bitmap[953] <= 1'b0;
		bitmap[954] <= 1'b0;
		bitmap[955] <= 1'b0;
		bitmap[956] <= 1'b0;
		bitmap[957] <= 1'b0;
		bitmap[958] <= 1'b0;
		bitmap[959] <= 1'b0;
		bitmap[960] <= 1'b0;
		bitmap[961] <= 1'b0;
		bitmap[962] <= 1'b0;
		bitmap[963] <= 1'b0;
		bitmap[964] <= 1'b0;
		bitmap[965] <= 1'b0;
		bitmap[966] <= 1'b0;
		bitmap[967] <= 1'b0;
		bitmap[968] <= 1'b0;
		bitmap[969] <= 1'b0;
		bitmap[970] <= 1'b0;
		bitmap[971] <= 1'b0;
		bitmap[972] <= 1'b0;
		bitmap[973] <= 1'b0;
		bitmap[974] <= 1'b0;
		bitmap[975] <= 1'b0;
		bitmap[976] <= 1'b0;
		bitmap[977] <= 1'b0;
		bitmap[978] <= 1'b0;
		bitmap[979] <= 1'b0;
		bitmap[980] <= 1'b0;
		bitmap[981] <= 1'b0;
		bitmap[982] <= 1'b0;
		bitmap[983] <= 1'b0;
		bitmap[984] <= 1'b0;
		bitmap[985] <= 1'b0;
		bitmap[986] <= 1'b0;
		bitmap[987] <= 1'b0;
		bitmap[988] <= 1'b0;
		bitmap[989] <= 1'b0;
		bitmap[990] <= 1'b0;
		bitmap[991] <= 1'b0;
		bitmap[992] <= 1'b0;
		bitmap[993] <= 1'b0;
		bitmap[994] <= 1'b0;
		bitmap[995] <= 1'b0;
		bitmap[996] <= 1'b0;
		bitmap[997] <= 1'b0;
		bitmap[998] <= 1'b0;
		bitmap[999] <= 1'b0;
		bitmap[1000] <= 1'b0;
		bitmap[1001] <= 1'b0;
		bitmap[1002] <= 1'b0;
		bitmap[1003] <= 1'b0;
		bitmap[1004] <= 1'b0;
		bitmap[1005] <= 1'b0;
		bitmap[1006] <= 1'b0;
		bitmap[1007] <= 1'b0;
		bitmap[1008] <= 1'b0;
		bitmap[1009] <= 1'b0;
		bitmap[1010] <= 1'b0;
		bitmap[1011] <= 1'b0;
		bitmap[1012] <= 1'b0;
		bitmap[1013] <= 1'b0;
		bitmap[1014] <= 1'b0;
		bitmap[1015] <= 1'b0;
		bitmap[1016] <= 1'b0;
		bitmap[1017] <= 1'b0;
		bitmap[1018] <= 1'b0;
		bitmap[1019] <= 1'b0;
		bitmap[1020] <= 1'b0;
		bitmap[1021] <= 1'b0;
		bitmap[1022] <= 1'b0;
		bitmap[1023] <= 1'b0;
		bitmap[1024] <= 1'b0;
		bitmap[1025] <= 1'b0;
		bitmap[1026] <= 1'b0;
		bitmap[1027] <= 1'b0;
		bitmap[1028] <= 1'b0;
		bitmap[1029] <= 1'b0;
		bitmap[1030] <= 1'b0;
		bitmap[1031] <= 1'b0;
		bitmap[1032] <= 1'b0;
		bitmap[1033] <= 1'b0;
		bitmap[1034] <= 1'b0;
		bitmap[1035] <= 1'b0;
		bitmap[1036] <= 1'b0;
		bitmap[1037] <= 1'b0;
		bitmap[1038] <= 1'b0;
		bitmap[1039] <= 1'b0;
		bitmap[1040] <= 1'b0;
		bitmap[1041] <= 1'b0;
		bitmap[1042] <= 1'b0;
		bitmap[1043] <= 1'b0;
		bitmap[1044] <= 1'b1;
		bitmap[1045] <= 1'b0;
		bitmap[1046] <= 1'b0;
		bitmap[1047] <= 1'b0;
		bitmap[1048] <= 1'b0;
		bitmap[1049] <= 1'b0;
		bitmap[1050] <= 1'b1;
		bitmap[1051] <= 1'b1;
		bitmap[1052] <= 1'b1;
		bitmap[1053] <= 1'b1;
		bitmap[1054] <= 1'b0;
		bitmap[1055] <= 1'b0;
		bitmap[1056] <= 1'b0;
		bitmap[1057] <= 1'b0;
		bitmap[1058] <= 1'b0;
		bitmap[1059] <= 1'b1;
		bitmap[1060] <= 1'b1;
		bitmap[1061] <= 1'b0;
		bitmap[1062] <= 1'b0;
		bitmap[1063] <= 1'b0;
		bitmap[1064] <= 1'b0;
		bitmap[1065] <= 1'b0;
		bitmap[1066] <= 1'b1;
		bitmap[1067] <= 1'b0;
		bitmap[1068] <= 1'b0;
		bitmap[1069] <= 1'b0;
		bitmap[1070] <= 1'b0;
		bitmap[1071] <= 1'b0;
		bitmap[1072] <= 1'b0;
		bitmap[1073] <= 1'b0;
		bitmap[1074] <= 1'b1;
		bitmap[1075] <= 1'b0;
		bitmap[1076] <= 1'b1;
		bitmap[1077] <= 1'b0;
		bitmap[1078] <= 1'b0;
		bitmap[1079] <= 1'b0;
		bitmap[1080] <= 1'b0;
		bitmap[1081] <= 1'b0;
		bitmap[1082] <= 1'b1;
		bitmap[1083] <= 1'b0;
		bitmap[1084] <= 1'b0;
		bitmap[1085] <= 1'b0;
		bitmap[1086] <= 1'b0;
		bitmap[1087] <= 1'b0;
		bitmap[1088] <= 1'b0;
		bitmap[1089] <= 1'b0;
		bitmap[1090] <= 1'b0;
		bitmap[1091] <= 1'b0;
		bitmap[1092] <= 1'b1;
		bitmap[1093] <= 1'b0;
		bitmap[1094] <= 1'b0;
		bitmap[1095] <= 1'b0;
		bitmap[1096] <= 1'b0;
		bitmap[1097] <= 1'b0;
		bitmap[1098] <= 1'b1;
		bitmap[1099] <= 1'b1;
		bitmap[1100] <= 1'b1;
		bitmap[1101] <= 1'b1;
		bitmap[1102] <= 1'b0;
		bitmap[1103] <= 1'b0;
		bitmap[1104] <= 1'b0;
		bitmap[1105] <= 1'b0;
		bitmap[1106] <= 1'b0;
		bitmap[1107] <= 1'b0;
		bitmap[1108] <= 1'b1;
		bitmap[1109] <= 1'b0;
		bitmap[1110] <= 1'b0;
		bitmap[1111] <= 1'b0;
		bitmap[1112] <= 1'b0;
		bitmap[1113] <= 1'b0;
		bitmap[1114] <= 1'b1;
		bitmap[1115] <= 1'b0;
		bitmap[1116] <= 1'b0;
		bitmap[1117] <= 1'b1;
		bitmap[1118] <= 1'b0;
		bitmap[1119] <= 1'b0;
		bitmap[1120] <= 1'b0;
		bitmap[1121] <= 1'b0;
		bitmap[1122] <= 1'b1;
		bitmap[1123] <= 1'b1;
		bitmap[1124] <= 1'b1;
		bitmap[1125] <= 1'b1;
		bitmap[1126] <= 1'b0;
		bitmap[1127] <= 1'b0;
		bitmap[1128] <= 1'b0;
		bitmap[1129] <= 1'b0;
		bitmap[1130] <= 1'b1;
		bitmap[1131] <= 1'b1;
		bitmap[1132] <= 1'b1;
		bitmap[1133] <= 1'b1;
		bitmap[1134] <= 1'b0;
		bitmap[1135] <= 1'b0;
		bitmap[1136] <= 1'b0;
		bitmap[1137] <= 1'b0;
		bitmap[1138] <= 1'b0;
		bitmap[1139] <= 1'b0;
		bitmap[1140] <= 1'b0;
		bitmap[1141] <= 1'b0;
		bitmap[1142] <= 1'b0;
		bitmap[1143] <= 1'b0;
		bitmap[1144] <= 1'b0;
		bitmap[1145] <= 1'b0;
		bitmap[1146] <= 1'b0;
		bitmap[1147] <= 1'b0;
		bitmap[1148] <= 1'b0;
		bitmap[1149] <= 1'b0;
		bitmap[1150] <= 1'b0;
		bitmap[1151] <= 1'b0;
		bitmap[1152] <= 1'b0;
		bitmap[1153] <= 1'b0;
		bitmap[1154] <= 1'b0;
		bitmap[1155] <= 1'b0;
		bitmap[1156] <= 1'b0;
		bitmap[1157] <= 1'b0;
		bitmap[1158] <= 1'b0;
		bitmap[1159] <= 1'b0;
		bitmap[1160] <= 1'b0;
		bitmap[1161] <= 1'b0;
		bitmap[1162] <= 1'b0;
		bitmap[1163] <= 1'b0;
		bitmap[1164] <= 1'b0;
		bitmap[1165] <= 1'b0;
		bitmap[1166] <= 1'b0;
		bitmap[1167] <= 1'b0;
		bitmap[1168] <= 1'b0;
		bitmap[1169] <= 1'b0;
		bitmap[1170] <= 1'b0;
		bitmap[1171] <= 1'b0;
		bitmap[1172] <= 1'b0;
		bitmap[1173] <= 1'b0;
		bitmap[1174] <= 1'b0;
		bitmap[1175] <= 1'b0;
		bitmap[1176] <= 1'b0;
		bitmap[1177] <= 1'b0;
		bitmap[1178] <= 1'b0;
		bitmap[1179] <= 1'b0;
		bitmap[1180] <= 1'b0;
		bitmap[1181] <= 1'b0;
		bitmap[1182] <= 1'b0;
		bitmap[1183] <= 1'b0;
		bitmap[1184] <= 1'b0;
		bitmap[1185] <= 1'b0;
		bitmap[1186] <= 1'b0;
		bitmap[1187] <= 1'b0;
		bitmap[1188] <= 1'b0;
		bitmap[1189] <= 1'b0;
		bitmap[1190] <= 1'b0;
		bitmap[1191] <= 1'b0;
		bitmap[1192] <= 1'b0;
		bitmap[1193] <= 1'b0;
		bitmap[1194] <= 1'b0;
		bitmap[1195] <= 1'b0;
		bitmap[1196] <= 1'b0;
		bitmap[1197] <= 1'b0;
		bitmap[1198] <= 1'b0;
		bitmap[1199] <= 1'b0;
		bitmap[1200] <= 1'b0;
		bitmap[1201] <= 1'b0;
		bitmap[1202] <= 1'b0;
		bitmap[1203] <= 1'b0;
		bitmap[1204] <= 1'b0;
		bitmap[1205] <= 1'b0;
		bitmap[1206] <= 1'b0;
		bitmap[1207] <= 1'b0;
		bitmap[1208] <= 1'b0;
		bitmap[1209] <= 1'b0;
		bitmap[1210] <= 1'b0;
		bitmap[1211] <= 1'b0;
		bitmap[1212] <= 1'b0;
		bitmap[1213] <= 1'b0;
		bitmap[1214] <= 1'b0;
		bitmap[1215] <= 1'b0;
		bitmap[1216] <= 1'b0;
		bitmap[1217] <= 1'b0;
		bitmap[1218] <= 1'b0;
		bitmap[1219] <= 1'b0;
		bitmap[1220] <= 1'b0;
		bitmap[1221] <= 1'b0;
		bitmap[1222] <= 1'b0;
		bitmap[1223] <= 1'b0;
		bitmap[1224] <= 1'b0;
		bitmap[1225] <= 1'b0;
		bitmap[1226] <= 1'b0;
		bitmap[1227] <= 1'b0;
		bitmap[1228] <= 1'b0;
		bitmap[1229] <= 1'b0;
		bitmap[1230] <= 1'b0;
		bitmap[1231] <= 1'b0;
		bitmap[1232] <= 1'b0;
		bitmap[1233] <= 1'b0;
		bitmap[1234] <= 1'b0;
		bitmap[1235] <= 1'b0;
		bitmap[1236] <= 1'b0;
		bitmap[1237] <= 1'b0;
		bitmap[1238] <= 1'b0;
		bitmap[1239] <= 1'b0;
		bitmap[1240] <= 1'b0;
		bitmap[1241] <= 1'b0;
		bitmap[1242] <= 1'b0;
		bitmap[1243] <= 1'b0;
		bitmap[1244] <= 1'b0;
		bitmap[1245] <= 1'b0;
		bitmap[1246] <= 1'b0;
		bitmap[1247] <= 1'b0;
		bitmap[1248] <= 1'b0;
		bitmap[1249] <= 1'b0;
		bitmap[1250] <= 1'b0;
		bitmap[1251] <= 1'b0;
		bitmap[1252] <= 1'b0;
		bitmap[1253] <= 1'b0;
		bitmap[1254] <= 1'b0;
		bitmap[1255] <= 1'b0;
		bitmap[1256] <= 1'b0;
		bitmap[1257] <= 1'b0;
		bitmap[1258] <= 1'b0;
		bitmap[1259] <= 1'b0;
		bitmap[1260] <= 1'b0;
		bitmap[1261] <= 1'b0;
		bitmap[1262] <= 1'b0;
		bitmap[1263] <= 1'b0;
		bitmap[1264] <= 1'b0;
		bitmap[1265] <= 1'b0;
		bitmap[1266] <= 1'b0;
		bitmap[1267] <= 1'b0;
		bitmap[1268] <= 1'b0;
		bitmap[1269] <= 1'b0;
		bitmap[1270] <= 1'b0;
		bitmap[1271] <= 1'b0;
		bitmap[1272] <= 1'b0;
		bitmap[1273] <= 1'b0;
		bitmap[1274] <= 1'b0;
		bitmap[1275] <= 1'b0;
		bitmap[1276] <= 1'b0;
		bitmap[1277] <= 1'b0;
		bitmap[1278] <= 1'b0;
		bitmap[1279] <= 1'b0;
		bitmap[1280] <= 1'b0;
		bitmap[1281] <= 1'b0;
		bitmap[1282] <= 1'b0;
		bitmap[1283] <= 1'b0;
		bitmap[1284] <= 1'b0;
		bitmap[1285] <= 1'b0;
		bitmap[1286] <= 1'b0;
		bitmap[1287] <= 1'b0;
		bitmap[1288] <= 1'b0;
		bitmap[1289] <= 1'b0;
		bitmap[1290] <= 1'b0;
		bitmap[1291] <= 1'b0;
		bitmap[1292] <= 1'b0;
		bitmap[1293] <= 1'b0;
		bitmap[1294] <= 1'b0;
		bitmap[1295] <= 1'b0;
		bitmap[1296] <= 1'b0;
		bitmap[1297] <= 1'b0;
		bitmap[1298] <= 1'b1;
		bitmap[1299] <= 1'b1;
		bitmap[1300] <= 1'b1;
		bitmap[1301] <= 1'b1;
		bitmap[1302] <= 1'b0;
		bitmap[1303] <= 1'b0;
		bitmap[1304] <= 1'b0;
		bitmap[1305] <= 1'b0;
		bitmap[1306] <= 1'b0;
		bitmap[1307] <= 1'b1;
		bitmap[1308] <= 1'b1;
		bitmap[1309] <= 1'b0;
		bitmap[1310] <= 1'b0;
		bitmap[1311] <= 1'b0;
		bitmap[1312] <= 1'b0;
		bitmap[1313] <= 1'b0;
		bitmap[1314] <= 1'b0;
		bitmap[1315] <= 1'b0;
		bitmap[1316] <= 1'b0;
		bitmap[1317] <= 1'b1;
		bitmap[1318] <= 1'b0;
		bitmap[1319] <= 1'b0;
		bitmap[1320] <= 1'b0;
		bitmap[1321] <= 1'b0;
		bitmap[1322] <= 1'b1;
		bitmap[1323] <= 1'b0;
		bitmap[1324] <= 1'b0;
		bitmap[1325] <= 1'b1;
		bitmap[1326] <= 1'b0;
		bitmap[1327] <= 1'b0;
		bitmap[1328] <= 1'b0;
		bitmap[1329] <= 1'b0;
		bitmap[1330] <= 1'b0;
		bitmap[1331] <= 1'b0;
		bitmap[1332] <= 1'b0;
		bitmap[1333] <= 1'b1;
		bitmap[1334] <= 1'b0;
		bitmap[1335] <= 1'b0;
		bitmap[1336] <= 1'b0;
		bitmap[1337] <= 1'b0;
		bitmap[1338] <= 1'b0;
		bitmap[1339] <= 1'b0;
		bitmap[1340] <= 1'b0;
		bitmap[1341] <= 1'b1;
		bitmap[1342] <= 1'b0;
		bitmap[1343] <= 1'b0;
		bitmap[1344] <= 1'b0;
		bitmap[1345] <= 1'b0;
		bitmap[1346] <= 1'b1;
		bitmap[1347] <= 1'b1;
		bitmap[1348] <= 1'b1;
		bitmap[1349] <= 1'b1;
		bitmap[1350] <= 1'b0;
		bitmap[1351] <= 1'b0;
		bitmap[1352] <= 1'b0;
		bitmap[1353] <= 1'b0;
		bitmap[1354] <= 1'b0;
		bitmap[1355] <= 1'b0;
		bitmap[1356] <= 1'b1;
		bitmap[1357] <= 1'b0;
		bitmap[1358] <= 1'b0;
		bitmap[1359] <= 1'b0;
		bitmap[1360] <= 1'b0;
		bitmap[1361] <= 1'b0;
		bitmap[1362] <= 1'b0;
		bitmap[1363] <= 1'b0;
		bitmap[1364] <= 1'b0;
		bitmap[1365] <= 1'b1;
		bitmap[1366] <= 1'b0;
		bitmap[1367] <= 1'b0;
		bitmap[1368] <= 1'b0;
		bitmap[1369] <= 1'b0;
		bitmap[1370] <= 1'b0;
		bitmap[1371] <= 1'b1;
		bitmap[1372] <= 1'b0;
		bitmap[1373] <= 1'b0;
		bitmap[1374] <= 1'b0;
		bitmap[1375] <= 1'b0;
		bitmap[1376] <= 1'b0;
		bitmap[1377] <= 1'b0;
		bitmap[1378] <= 1'b1;
		bitmap[1379] <= 1'b1;
		bitmap[1380] <= 1'b1;
		bitmap[1381] <= 1'b1;
		bitmap[1382] <= 1'b0;
		bitmap[1383] <= 1'b0;
		bitmap[1384] <= 1'b0;
		bitmap[1385] <= 1'b0;
		bitmap[1386] <= 1'b1;
		bitmap[1387] <= 1'b1;
		bitmap[1388] <= 1'b1;
		bitmap[1389] <= 1'b1;
		bitmap[1390] <= 1'b0;
		bitmap[1391] <= 1'b0;
		bitmap[1392] <= 1'b0;
		bitmap[1393] <= 1'b0;
		bitmap[1394] <= 1'b0;
		bitmap[1395] <= 1'b0;
		bitmap[1396] <= 1'b0;
		bitmap[1397] <= 1'b0;
		bitmap[1398] <= 1'b0;
		bitmap[1399] <= 1'b0;
		bitmap[1400] <= 1'b0;
		bitmap[1401] <= 1'b0;
		bitmap[1402] <= 1'b0;
		bitmap[1403] <= 1'b0;
		bitmap[1404] <= 1'b0;
		bitmap[1405] <= 1'b0;
		bitmap[1406] <= 1'b0;
		bitmap[1407] <= 1'b0;
		bitmap[1408] <= 1'b0;
		bitmap[1409] <= 1'b0;
		bitmap[1410] <= 1'b0;
		bitmap[1411] <= 1'b0;
		bitmap[1412] <= 1'b0;
		bitmap[1413] <= 1'b0;
		bitmap[1414] <= 1'b0;
		bitmap[1415] <= 1'b0;
		bitmap[1416] <= 1'b0;
		bitmap[1417] <= 1'b0;
		bitmap[1418] <= 1'b0;
		bitmap[1419] <= 1'b0;
		bitmap[1420] <= 1'b0;
		bitmap[1421] <= 1'b0;
		bitmap[1422] <= 1'b0;
		bitmap[1423] <= 1'b0;
		bitmap[1424] <= 1'b0;
		bitmap[1425] <= 1'b0;
		bitmap[1426] <= 1'b0;
		bitmap[1427] <= 1'b0;
		bitmap[1428] <= 1'b0;
		bitmap[1429] <= 1'b0;
		bitmap[1430] <= 1'b0;
		bitmap[1431] <= 1'b0;
		bitmap[1432] <= 1'b0;
		bitmap[1433] <= 1'b0;
		bitmap[1434] <= 1'b0;
		bitmap[1435] <= 1'b0;
		bitmap[1436] <= 1'b0;
		bitmap[1437] <= 1'b0;
		bitmap[1438] <= 1'b0;
		bitmap[1439] <= 1'b0;
		bitmap[1440] <= 1'b0;
		bitmap[1441] <= 1'b0;
		bitmap[1442] <= 1'b0;
		bitmap[1443] <= 1'b0;
		bitmap[1444] <= 1'b0;
		bitmap[1445] <= 1'b0;
		bitmap[1446] <= 1'b0;
		bitmap[1447] <= 1'b0;
		bitmap[1448] <= 1'b0;
		bitmap[1449] <= 1'b0;
		bitmap[1450] <= 1'b0;
		bitmap[1451] <= 1'b0;
		bitmap[1452] <= 1'b0;
		bitmap[1453] <= 1'b0;
		bitmap[1454] <= 1'b0;
		bitmap[1455] <= 1'b0;
		bitmap[1456] <= 1'b0;
		bitmap[1457] <= 1'b0;
		bitmap[1458] <= 1'b0;
		bitmap[1459] <= 1'b0;
		bitmap[1460] <= 1'b0;
		bitmap[1461] <= 1'b0;
		bitmap[1462] <= 1'b0;
		bitmap[1463] <= 1'b0;
		bitmap[1464] <= 1'b0;
		bitmap[1465] <= 1'b0;
		bitmap[1466] <= 1'b0;
		bitmap[1467] <= 1'b0;
		bitmap[1468] <= 1'b0;
		bitmap[1469] <= 1'b0;
		bitmap[1470] <= 1'b0;
		bitmap[1471] <= 1'b0;
		bitmap[1472] <= 1'b0;
		bitmap[1473] <= 1'b0;
		bitmap[1474] <= 1'b0;
		bitmap[1475] <= 1'b0;
		bitmap[1476] <= 1'b0;
		bitmap[1477] <= 1'b0;
		bitmap[1478] <= 1'b0;
		bitmap[1479] <= 1'b0;
		bitmap[1480] <= 1'b0;
		bitmap[1481] <= 1'b0;
		bitmap[1482] <= 1'b0;
		bitmap[1483] <= 1'b0;
		bitmap[1484] <= 1'b0;
		bitmap[1485] <= 1'b0;
		bitmap[1486] <= 1'b0;
		bitmap[1487] <= 1'b0;
		bitmap[1488] <= 1'b0;
		bitmap[1489] <= 1'b0;
		bitmap[1490] <= 1'b0;
		bitmap[1491] <= 1'b0;
		bitmap[1492] <= 1'b0;
		bitmap[1493] <= 1'b0;
		bitmap[1494] <= 1'b0;
		bitmap[1495] <= 1'b0;
		bitmap[1496] <= 1'b0;
		bitmap[1497] <= 1'b0;
		bitmap[1498] <= 1'b0;
		bitmap[1499] <= 1'b0;
		bitmap[1500] <= 1'b0;
		bitmap[1501] <= 1'b0;
		bitmap[1502] <= 1'b0;
		bitmap[1503] <= 1'b0;
		bitmap[1504] <= 1'b0;
		bitmap[1505] <= 1'b0;
		bitmap[1506] <= 1'b0;
		bitmap[1507] <= 1'b0;
		bitmap[1508] <= 1'b0;
		bitmap[1509] <= 1'b0;
		bitmap[1510] <= 1'b0;
		bitmap[1511] <= 1'b0;
		bitmap[1512] <= 1'b0;
		bitmap[1513] <= 1'b0;
		bitmap[1514] <= 1'b0;
		bitmap[1515] <= 1'b0;
		bitmap[1516] <= 1'b0;
		bitmap[1517] <= 1'b0;
		bitmap[1518] <= 1'b0;
		bitmap[1519] <= 1'b0;
		bitmap[1520] <= 1'b0;
		bitmap[1521] <= 1'b0;
		bitmap[1522] <= 1'b0;
		bitmap[1523] <= 1'b0;
		bitmap[1524] <= 1'b0;
		bitmap[1525] <= 1'b0;
		bitmap[1526] <= 1'b0;
		bitmap[1527] <= 1'b0;
		bitmap[1528] <= 1'b0;
		bitmap[1529] <= 1'b0;
		bitmap[1530] <= 1'b0;
		bitmap[1531] <= 1'b0;
		bitmap[1532] <= 1'b0;
		bitmap[1533] <= 1'b0;
		bitmap[1534] <= 1'b0;
		bitmap[1535] <= 1'b0;
		bitmap[1536] <= 1'b0;
		bitmap[1537] <= 1'b0;
		bitmap[1538] <= 1'b0;
		bitmap[1539] <= 1'b0;
		bitmap[1540] <= 1'b0;
		bitmap[1541] <= 1'b0;
		bitmap[1542] <= 1'b0;
		bitmap[1543] <= 1'b0;
		bitmap[1544] <= 1'b0;
		bitmap[1545] <= 1'b0;
		bitmap[1546] <= 1'b0;
		bitmap[1547] <= 1'b0;
		bitmap[1548] <= 1'b0;
		bitmap[1549] <= 1'b0;
		bitmap[1550] <= 1'b0;
		bitmap[1551] <= 1'b0;
		bitmap[1552] <= 1'b0;
		bitmap[1553] <= 1'b0;
		bitmap[1554] <= 1'b1;
		bitmap[1555] <= 1'b1;
		bitmap[1556] <= 1'b1;
		bitmap[1557] <= 1'b1;
		bitmap[1558] <= 1'b0;
		bitmap[1559] <= 1'b0;
		bitmap[1560] <= 1'b0;
		bitmap[1561] <= 1'b0;
		bitmap[1562] <= 1'b0;
		bitmap[1563] <= 1'b0;
		bitmap[1564] <= 1'b1;
		bitmap[1565] <= 1'b1;
		bitmap[1566] <= 1'b0;
		bitmap[1567] <= 1'b0;
		bitmap[1568] <= 1'b0;
		bitmap[1569] <= 1'b0;
		bitmap[1570] <= 1'b1;
		bitmap[1571] <= 1'b0;
		bitmap[1572] <= 1'b0;
		bitmap[1573] <= 1'b0;
		bitmap[1574] <= 1'b0;
		bitmap[1575] <= 1'b0;
		bitmap[1576] <= 1'b0;
		bitmap[1577] <= 1'b0;
		bitmap[1578] <= 1'b0;
		bitmap[1579] <= 1'b1;
		bitmap[1580] <= 1'b0;
		bitmap[1581] <= 1'b1;
		bitmap[1582] <= 1'b0;
		bitmap[1583] <= 1'b0;
		bitmap[1584] <= 1'b0;
		bitmap[1585] <= 1'b0;
		bitmap[1586] <= 1'b1;
		bitmap[1587] <= 1'b0;
		bitmap[1588] <= 1'b0;
		bitmap[1589] <= 1'b0;
		bitmap[1590] <= 1'b0;
		bitmap[1591] <= 1'b0;
		bitmap[1592] <= 1'b0;
		bitmap[1593] <= 1'b0;
		bitmap[1594] <= 1'b1;
		bitmap[1595] <= 1'b0;
		bitmap[1596] <= 1'b0;
		bitmap[1597] <= 1'b1;
		bitmap[1598] <= 1'b0;
		bitmap[1599] <= 1'b0;
		bitmap[1600] <= 1'b0;
		bitmap[1601] <= 1'b0;
		bitmap[1602] <= 1'b1;
		bitmap[1603] <= 1'b1;
		bitmap[1604] <= 1'b1;
		bitmap[1605] <= 1'b1;
		bitmap[1606] <= 1'b0;
		bitmap[1607] <= 1'b0;
		bitmap[1608] <= 1'b0;
		bitmap[1609] <= 1'b0;
		bitmap[1610] <= 1'b1;
		bitmap[1611] <= 1'b1;
		bitmap[1612] <= 1'b1;
		bitmap[1613] <= 1'b1;
		bitmap[1614] <= 1'b1;
		bitmap[1615] <= 1'b0;
		bitmap[1616] <= 1'b0;
		bitmap[1617] <= 1'b0;
		bitmap[1618] <= 1'b1;
		bitmap[1619] <= 1'b0;
		bitmap[1620] <= 1'b0;
		bitmap[1621] <= 1'b1;
		bitmap[1622] <= 1'b0;
		bitmap[1623] <= 1'b0;
		bitmap[1624] <= 1'b0;
		bitmap[1625] <= 1'b0;
		bitmap[1626] <= 1'b0;
		bitmap[1627] <= 1'b0;
		bitmap[1628] <= 1'b0;
		bitmap[1629] <= 1'b1;
		bitmap[1630] <= 1'b0;
		bitmap[1631] <= 1'b0;
		bitmap[1632] <= 1'b0;
		bitmap[1633] <= 1'b0;
		bitmap[1634] <= 1'b1;
		bitmap[1635] <= 1'b1;
		bitmap[1636] <= 1'b1;
		bitmap[1637] <= 1'b1;
		bitmap[1638] <= 1'b0;
		bitmap[1639] <= 1'b0;
		bitmap[1640] <= 1'b0;
		bitmap[1641] <= 1'b0;
		bitmap[1642] <= 1'b0;
		bitmap[1643] <= 1'b0;
		bitmap[1644] <= 1'b0;
		bitmap[1645] <= 1'b1;
		bitmap[1646] <= 1'b0;
		bitmap[1647] <= 1'b0;
		bitmap[1648] <= 1'b0;
		bitmap[1649] <= 1'b0;
		bitmap[1650] <= 1'b0;
		bitmap[1651] <= 1'b0;
		bitmap[1652] <= 1'b0;
		bitmap[1653] <= 1'b0;
		bitmap[1654] <= 1'b0;
		bitmap[1655] <= 1'b0;
		bitmap[1656] <= 1'b0;
		bitmap[1657] <= 1'b0;
		bitmap[1658] <= 1'b0;
		bitmap[1659] <= 1'b0;
		bitmap[1660] <= 1'b0;
		bitmap[1661] <= 1'b0;
		bitmap[1662] <= 1'b0;
		bitmap[1663] <= 1'b0;
		bitmap[1664] <= 1'b0;
		bitmap[1665] <= 1'b0;
		bitmap[1666] <= 1'b0;
		bitmap[1667] <= 1'b0;
		bitmap[1668] <= 1'b0;
		bitmap[1669] <= 1'b0;
		bitmap[1670] <= 1'b0;
		bitmap[1671] <= 1'b0;
		bitmap[1672] <= 1'b0;
		bitmap[1673] <= 1'b0;
		bitmap[1674] <= 1'b0;
		bitmap[1675] <= 1'b0;
		bitmap[1676] <= 1'b0;
		bitmap[1677] <= 1'b0;
		bitmap[1678] <= 1'b0;
		bitmap[1679] <= 1'b0;
		bitmap[1680] <= 1'b0;
		bitmap[1681] <= 1'b0;
		bitmap[1682] <= 1'b0;
		bitmap[1683] <= 1'b0;
		bitmap[1684] <= 1'b0;
		bitmap[1685] <= 1'b0;
		bitmap[1686] <= 1'b0;
		bitmap[1687] <= 1'b0;
		bitmap[1688] <= 1'b0;
		bitmap[1689] <= 1'b0;
		bitmap[1690] <= 1'b0;
		bitmap[1691] <= 1'b0;
		bitmap[1692] <= 1'b0;
		bitmap[1693] <= 1'b0;
		bitmap[1694] <= 1'b0;
		bitmap[1695] <= 1'b0;
		bitmap[1696] <= 1'b0;
		bitmap[1697] <= 1'b0;
		bitmap[1698] <= 1'b0;
		bitmap[1699] <= 1'b0;
		bitmap[1700] <= 1'b0;
		bitmap[1701] <= 1'b0;
		bitmap[1702] <= 1'b0;
		bitmap[1703] <= 1'b0;
		bitmap[1704] <= 1'b0;
		bitmap[1705] <= 1'b0;
		bitmap[1706] <= 1'b0;
		bitmap[1707] <= 1'b0;
		bitmap[1708] <= 1'b0;
		bitmap[1709] <= 1'b0;
		bitmap[1710] <= 1'b0;
		bitmap[1711] <= 1'b0;
		bitmap[1712] <= 1'b0;
		bitmap[1713] <= 1'b0;
		bitmap[1714] <= 1'b0;
		bitmap[1715] <= 1'b0;
		bitmap[1716] <= 1'b0;
		bitmap[1717] <= 1'b0;
		bitmap[1718] <= 1'b0;
		bitmap[1719] <= 1'b0;
		bitmap[1720] <= 1'b0;
		bitmap[1721] <= 1'b0;
		bitmap[1722] <= 1'b0;
		bitmap[1723] <= 1'b0;
		bitmap[1724] <= 1'b0;
		bitmap[1725] <= 1'b0;
		bitmap[1726] <= 1'b0;
		bitmap[1727] <= 1'b0;
		bitmap[1728] <= 1'b0;
		bitmap[1729] <= 1'b0;
		bitmap[1730] <= 1'b0;
		bitmap[1731] <= 1'b0;
		bitmap[1732] <= 1'b0;
		bitmap[1733] <= 1'b0;
		bitmap[1734] <= 1'b0;
		bitmap[1735] <= 1'b0;
		bitmap[1736] <= 1'b0;
		bitmap[1737] <= 1'b0;
		bitmap[1738] <= 1'b0;
		bitmap[1739] <= 1'b0;
		bitmap[1740] <= 1'b0;
		bitmap[1741] <= 1'b0;
		bitmap[1742] <= 1'b0;
		bitmap[1743] <= 1'b0;
		bitmap[1744] <= 1'b0;
		bitmap[1745] <= 1'b0;
		bitmap[1746] <= 1'b0;
		bitmap[1747] <= 1'b0;
		bitmap[1748] <= 1'b0;
		bitmap[1749] <= 1'b0;
		bitmap[1750] <= 1'b0;
		bitmap[1751] <= 1'b0;
		bitmap[1752] <= 1'b0;
		bitmap[1753] <= 1'b0;
		bitmap[1754] <= 1'b0;
		bitmap[1755] <= 1'b0;
		bitmap[1756] <= 1'b0;
		bitmap[1757] <= 1'b0;
		bitmap[1758] <= 1'b0;
		bitmap[1759] <= 1'b0;
		bitmap[1760] <= 1'b0;
		bitmap[1761] <= 1'b0;
		bitmap[1762] <= 1'b0;
		bitmap[1763] <= 1'b0;
		bitmap[1764] <= 1'b0;
		bitmap[1765] <= 1'b0;
		bitmap[1766] <= 1'b0;
		bitmap[1767] <= 1'b0;
		bitmap[1768] <= 1'b0;
		bitmap[1769] <= 1'b0;
		bitmap[1770] <= 1'b0;
		bitmap[1771] <= 1'b0;
		bitmap[1772] <= 1'b0;
		bitmap[1773] <= 1'b0;
		bitmap[1774] <= 1'b0;
		bitmap[1775] <= 1'b0;
		bitmap[1776] <= 1'b0;
		bitmap[1777] <= 1'b0;
		bitmap[1778] <= 1'b0;
		bitmap[1779] <= 1'b0;
		bitmap[1780] <= 1'b0;
		bitmap[1781] <= 1'b0;
		bitmap[1782] <= 1'b0;
		bitmap[1783] <= 1'b0;
		bitmap[1784] <= 1'b0;
		bitmap[1785] <= 1'b0;
		bitmap[1786] <= 1'b0;
		bitmap[1787] <= 1'b0;
		bitmap[1788] <= 1'b0;
		bitmap[1789] <= 1'b0;
		bitmap[1790] <= 1'b0;
		bitmap[1791] <= 1'b0;
		bitmap[1792] <= 1'b0;
		bitmap[1793] <= 1'b0;
		bitmap[1794] <= 1'b0;
		bitmap[1795] <= 1'b0;
		bitmap[1796] <= 1'b0;
		bitmap[1797] <= 1'b0;
		bitmap[1798] <= 1'b0;
		bitmap[1799] <= 1'b0;
		bitmap[1800] <= 1'b0;
		bitmap[1801] <= 1'b0;
		bitmap[1802] <= 1'b0;
		bitmap[1803] <= 1'b0;
		bitmap[1804] <= 1'b0;
		bitmap[1805] <= 1'b0;
		bitmap[1806] <= 1'b0;
		bitmap[1807] <= 1'b0;
		bitmap[1808] <= 1'b0;
		bitmap[1809] <= 1'b0;
		bitmap[1810] <= 1'b0;
		bitmap[1811] <= 1'b0;
		bitmap[1812] <= 1'b1;
		bitmap[1813] <= 1'b0;
		bitmap[1814] <= 1'b0;
		bitmap[1815] <= 1'b0;
		bitmap[1816] <= 1'b0;
		bitmap[1817] <= 1'b0;
		bitmap[1818] <= 1'b0;
		bitmap[1819] <= 1'b1;
		bitmap[1820] <= 1'b1;
		bitmap[1821] <= 1'b0;
		bitmap[1822] <= 1'b0;
		bitmap[1823] <= 1'b0;
		bitmap[1824] <= 1'b0;
		bitmap[1825] <= 1'b0;
		bitmap[1826] <= 1'b0;
		bitmap[1827] <= 1'b1;
		bitmap[1828] <= 1'b1;
		bitmap[1829] <= 1'b0;
		bitmap[1830] <= 1'b0;
		bitmap[1831] <= 1'b0;
		bitmap[1832] <= 1'b0;
		bitmap[1833] <= 1'b0;
		bitmap[1834] <= 1'b1;
		bitmap[1835] <= 1'b0;
		bitmap[1836] <= 1'b0;
		bitmap[1837] <= 1'b1;
		bitmap[1838] <= 1'b0;
		bitmap[1839] <= 1'b0;
		bitmap[1840] <= 1'b0;
		bitmap[1841] <= 1'b0;
		bitmap[1842] <= 1'b1;
		bitmap[1843] <= 1'b0;
		bitmap[1844] <= 1'b1;
		bitmap[1845] <= 1'b0;
		bitmap[1846] <= 1'b0;
		bitmap[1847] <= 1'b0;
		bitmap[1848] <= 1'b0;
		bitmap[1849] <= 1'b0;
		bitmap[1850] <= 1'b0;
		bitmap[1851] <= 1'b0;
		bitmap[1852] <= 1'b0;
		bitmap[1853] <= 1'b1;
		bitmap[1854] <= 1'b0;
		bitmap[1855] <= 1'b0;
		bitmap[1856] <= 1'b0;
		bitmap[1857] <= 1'b0;
		bitmap[1858] <= 1'b0;
		bitmap[1859] <= 1'b0;
		bitmap[1860] <= 1'b1;
		bitmap[1861] <= 1'b0;
		bitmap[1862] <= 1'b0;
		bitmap[1863] <= 1'b0;
		bitmap[1864] <= 1'b0;
		bitmap[1865] <= 1'b0;
		bitmap[1866] <= 1'b0;
		bitmap[1867] <= 1'b0;
		bitmap[1868] <= 1'b1;
		bitmap[1869] <= 1'b0;
		bitmap[1870] <= 1'b0;
		bitmap[1871] <= 1'b0;
		bitmap[1872] <= 1'b0;
		bitmap[1873] <= 1'b0;
		bitmap[1874] <= 1'b0;
		bitmap[1875] <= 1'b0;
		bitmap[1876] <= 1'b1;
		bitmap[1877] <= 1'b0;
		bitmap[1878] <= 1'b0;
		bitmap[1879] <= 1'b0;
		bitmap[1880] <= 1'b0;
		bitmap[1881] <= 1'b0;
		bitmap[1882] <= 1'b0;
		bitmap[1883] <= 1'b1;
		bitmap[1884] <= 1'b0;
		bitmap[1885] <= 1'b0;
		bitmap[1886] <= 1'b0;
		bitmap[1887] <= 1'b0;
		bitmap[1888] <= 1'b0;
		bitmap[1889] <= 1'b0;
		bitmap[1890] <= 1'b1;
		bitmap[1891] <= 1'b1;
		bitmap[1892] <= 1'b1;
		bitmap[1893] <= 1'b1;
		bitmap[1894] <= 1'b0;
		bitmap[1895] <= 1'b0;
		bitmap[1896] <= 1'b0;
		bitmap[1897] <= 1'b0;
		bitmap[1898] <= 1'b1;
		bitmap[1899] <= 1'b1;
		bitmap[1900] <= 1'b1;
		bitmap[1901] <= 1'b1;
		bitmap[1902] <= 1'b0;
		bitmap[1903] <= 1'b0;
		bitmap[1904] <= 1'b0;
		bitmap[1905] <= 1'b0;
		bitmap[1906] <= 1'b0;
		bitmap[1907] <= 1'b0;
		bitmap[1908] <= 1'b0;
		bitmap[1909] <= 1'b0;
		bitmap[1910] <= 1'b0;
		bitmap[1911] <= 1'b0;
		bitmap[1912] <= 1'b0;
		bitmap[1913] <= 1'b0;
		bitmap[1914] <= 1'b0;
		bitmap[1915] <= 1'b0;
		bitmap[1916] <= 1'b0;
		bitmap[1917] <= 1'b0;
		bitmap[1918] <= 1'b0;
		bitmap[1919] <= 1'b0;
		bitmap[1920] <= 1'b0;
		bitmap[1921] <= 1'b0;
		bitmap[1922] <= 1'b0;
		bitmap[1923] <= 1'b0;
		bitmap[1924] <= 1'b0;
		bitmap[1925] <= 1'b0;
		bitmap[1926] <= 1'b0;
		bitmap[1927] <= 1'b0;
		bitmap[1928] <= 1'b0;
		bitmap[1929] <= 1'b0;
		bitmap[1930] <= 1'b0;
		bitmap[1931] <= 1'b0;
		bitmap[1932] <= 1'b0;
		bitmap[1933] <= 1'b0;
		bitmap[1934] <= 1'b0;
		bitmap[1935] <= 1'b0;
		bitmap[1936] <= 1'b0;
		bitmap[1937] <= 1'b0;
		bitmap[1938] <= 1'b1;
		bitmap[1939] <= 1'b1;
		bitmap[1940] <= 1'b1;
		bitmap[1941] <= 1'b1;
		bitmap[1942] <= 1'b0;
		bitmap[1943] <= 1'b0;
		bitmap[1944] <= 1'b0;
		bitmap[1945] <= 1'b0;
		bitmap[1946] <= 1'b0;
		bitmap[1947] <= 1'b0;
		bitmap[1948] <= 1'b0;
		bitmap[1949] <= 1'b0;
		bitmap[1950] <= 1'b0;
		bitmap[1951] <= 1'b0;
		bitmap[1952] <= 1'b0;
		bitmap[1953] <= 1'b0;
		bitmap[1954] <= 1'b1;
		bitmap[1955] <= 1'b0;
		bitmap[1956] <= 1'b0;
		bitmap[1957] <= 1'b1;
		bitmap[1958] <= 1'b0;
		bitmap[1959] <= 1'b0;
		bitmap[1960] <= 1'b0;
		bitmap[1961] <= 1'b0;
		bitmap[1962] <= 1'b0;
		bitmap[1963] <= 1'b0;
		bitmap[1964] <= 1'b0;
		bitmap[1965] <= 1'b0;
		bitmap[1966] <= 1'b0;
		bitmap[1967] <= 1'b0;
		bitmap[1968] <= 1'b0;
		bitmap[1969] <= 1'b0;
		bitmap[1970] <= 1'b1;
		bitmap[1971] <= 1'b0;
		bitmap[1972] <= 1'b0;
		bitmap[1973] <= 1'b1;
		bitmap[1974] <= 1'b0;
		bitmap[1975] <= 1'b0;
		bitmap[1976] <= 1'b0;
		bitmap[1977] <= 1'b0;
		bitmap[1978] <= 1'b0;
		bitmap[1979] <= 1'b0;
		bitmap[1980] <= 1'b0;
		bitmap[1981] <= 1'b0;
		bitmap[1982] <= 1'b0;
		bitmap[1983] <= 1'b0;
		bitmap[1984] <= 1'b0;
		bitmap[1985] <= 1'b0;
		bitmap[1986] <= 1'b1;
		bitmap[1987] <= 1'b1;
		bitmap[1988] <= 1'b1;
		bitmap[1989] <= 1'b1;
		bitmap[1990] <= 1'b0;
		bitmap[1991] <= 1'b0;
		bitmap[1992] <= 1'b0;
		bitmap[1993] <= 1'b0;
		bitmap[1994] <= 1'b0;
		bitmap[1995] <= 1'b0;
		bitmap[1996] <= 1'b0;
		bitmap[1997] <= 1'b0;
		bitmap[1998] <= 1'b0;
		bitmap[1999] <= 1'b0;
		bitmap[2000] <= 1'b0;
		bitmap[2001] <= 1'b0;
		bitmap[2002] <= 1'b1;
		bitmap[2003] <= 1'b0;
		bitmap[2004] <= 1'b0;
		bitmap[2005] <= 1'b1;
		bitmap[2006] <= 1'b0;
		bitmap[2007] <= 1'b0;
		bitmap[2008] <= 1'b0;
		bitmap[2009] <= 1'b0;
		bitmap[2010] <= 1'b0;
		bitmap[2011] <= 1'b0;
		bitmap[2012] <= 1'b0;
		bitmap[2013] <= 1'b0;
		bitmap[2014] <= 1'b0;
		bitmap[2015] <= 1'b0;
		bitmap[2016] <= 1'b0;
		bitmap[2017] <= 1'b0;
		bitmap[2018] <= 1'b1;
		bitmap[2019] <= 1'b1;
		bitmap[2020] <= 1'b1;
		bitmap[2021] <= 1'b1;
		bitmap[2022] <= 1'b0;
		bitmap[2023] <= 1'b0;
		bitmap[2024] <= 1'b0;
		bitmap[2025] <= 1'b0;
		bitmap[2026] <= 1'b0;
		bitmap[2027] <= 1'b0;
		bitmap[2028] <= 1'b0;
		bitmap[2029] <= 1'b0;
		bitmap[2030] <= 1'b0;
		bitmap[2031] <= 1'b0;
		bitmap[2032] <= 1'b0;
		bitmap[2033] <= 1'b0;
		bitmap[2034] <= 1'b0;
		bitmap[2035] <= 1'b0;
		bitmap[2036] <= 1'b0;
		bitmap[2037] <= 1'b0;
		bitmap[2038] <= 1'b0;
		bitmap[2039] <= 1'b0;
		bitmap[2040] <= 1'b0;
		bitmap[2041] <= 1'b0;
		bitmap[2042] <= 1'b0;
		bitmap[2043] <= 1'b0;
		bitmap[2044] <= 1'b0;
		bitmap[2045] <= 1'b0;
		bitmap[2046] <= 1'b0;
		bitmap[2047] <= 1'b0;
		bitmap[2048] <= 1'b0;
		bitmap[2049] <= 1'b0;
		bitmap[2050] <= 1'b0;
		bitmap[2051] <= 1'b0;
		bitmap[2052] <= 1'b0;
		bitmap[2053] <= 1'b0;
		bitmap[2054] <= 1'b0;
		bitmap[2055] <= 1'b0;
		bitmap[2056] <= 1'b0;
		bitmap[2057] <= 1'b0;
		bitmap[2058] <= 1'b0;
		bitmap[2059] <= 1'b0;
		bitmap[2060] <= 1'b0;
		bitmap[2061] <= 1'b0;
		bitmap[2062] <= 1'b0;
		bitmap[2063] <= 1'b0;
		bitmap[2064] <= 1'b0;
		bitmap[2065] <= 1'b0;
		bitmap[2066] <= 1'b0;
		bitmap[2067] <= 1'b1;
		bitmap[2068] <= 1'b1;
		bitmap[2069] <= 1'b0;
		bitmap[2070] <= 1'b0;
		bitmap[2071] <= 1'b0;
		bitmap[2072] <= 1'b0;
		bitmap[2073] <= 1'b0;
		bitmap[2074] <= 1'b1;
		bitmap[2075] <= 1'b1;
		bitmap[2076] <= 1'b1;
		bitmap[2077] <= 1'b1;
		bitmap[2078] <= 1'b0;
		bitmap[2079] <= 1'b0;
		bitmap[2080] <= 1'b0;
		bitmap[2081] <= 1'b0;
		bitmap[2082] <= 1'b1;
		bitmap[2083] <= 1'b0;
		bitmap[2084] <= 1'b0;
		bitmap[2085] <= 1'b1;
		bitmap[2086] <= 1'b0;
		bitmap[2087] <= 1'b0;
		bitmap[2088] <= 1'b0;
		bitmap[2089] <= 1'b0;
		bitmap[2090] <= 1'b1;
		bitmap[2091] <= 1'b0;
		bitmap[2092] <= 1'b0;
		bitmap[2093] <= 1'b0;
		bitmap[2094] <= 1'b0;
		bitmap[2095] <= 1'b0;
		bitmap[2096] <= 1'b0;
		bitmap[2097] <= 1'b0;
		bitmap[2098] <= 1'b0;
		bitmap[2099] <= 1'b0;
		bitmap[2100] <= 1'b0;
		bitmap[2101] <= 1'b1;
		bitmap[2102] <= 1'b0;
		bitmap[2103] <= 1'b0;
		bitmap[2104] <= 1'b0;
		bitmap[2105] <= 1'b0;
		bitmap[2106] <= 1'b1;
		bitmap[2107] <= 1'b0;
		bitmap[2108] <= 1'b0;
		bitmap[2109] <= 1'b0;
		bitmap[2110] <= 1'b0;
		bitmap[2111] <= 1'b0;
		bitmap[2112] <= 1'b0;
		bitmap[2113] <= 1'b0;
		bitmap[2114] <= 1'b0;
		bitmap[2115] <= 1'b0;
		bitmap[2116] <= 1'b1;
		bitmap[2117] <= 1'b0;
		bitmap[2118] <= 1'b0;
		bitmap[2119] <= 1'b0;
		bitmap[2120] <= 1'b0;
		bitmap[2121] <= 1'b0;
		bitmap[2122] <= 1'b1;
		bitmap[2123] <= 1'b1;
		bitmap[2124] <= 1'b1;
		bitmap[2125] <= 1'b1;
		bitmap[2126] <= 1'b0;
		bitmap[2127] <= 1'b0;
		bitmap[2128] <= 1'b0;
		bitmap[2129] <= 1'b0;
		bitmap[2130] <= 1'b0;
		bitmap[2131] <= 1'b1;
		bitmap[2132] <= 1'b0;
		bitmap[2133] <= 1'b0;
		bitmap[2134] <= 1'b0;
		bitmap[2135] <= 1'b0;
		bitmap[2136] <= 1'b0;
		bitmap[2137] <= 1'b0;
		bitmap[2138] <= 1'b0;
		bitmap[2139] <= 1'b0;
		bitmap[2140] <= 1'b0;
		bitmap[2141] <= 1'b1;
		bitmap[2142] <= 1'b0;
		bitmap[2143] <= 1'b0;
		bitmap[2144] <= 1'b0;
		bitmap[2145] <= 1'b0;
		bitmap[2146] <= 1'b1;
		bitmap[2147] <= 1'b1;
		bitmap[2148] <= 1'b1;
		bitmap[2149] <= 1'b1;
		bitmap[2150] <= 1'b0;
		bitmap[2151] <= 1'b0;
		bitmap[2152] <= 1'b0;
		bitmap[2153] <= 1'b0;
		bitmap[2154] <= 1'b1;
		bitmap[2155] <= 1'b1;
		bitmap[2156] <= 1'b1;
		bitmap[2157] <= 1'b1;
		bitmap[2158] <= 1'b0;
		bitmap[2159] <= 1'b0;
		bitmap[2160] <= 1'b0;
		bitmap[2161] <= 1'b0;
		bitmap[2162] <= 1'b0;
		bitmap[2163] <= 1'b0;
		bitmap[2164] <= 1'b0;
		bitmap[2165] <= 1'b0;
		bitmap[2166] <= 1'b0;
		bitmap[2167] <= 1'b0;
		bitmap[2168] <= 1'b0;
		bitmap[2169] <= 1'b0;
		bitmap[2170] <= 1'b0;
		bitmap[2171] <= 1'b0;
		bitmap[2172] <= 1'b0;
		bitmap[2173] <= 1'b0;
		bitmap[2174] <= 1'b0;
		bitmap[2175] <= 1'b0;
		bitmap[2176] <= 1'b0;
		bitmap[2177] <= 1'b0;
		bitmap[2178] <= 1'b0;
		bitmap[2179] <= 1'b0;
		bitmap[2180] <= 1'b0;
		bitmap[2181] <= 1'b0;
		bitmap[2182] <= 1'b0;
		bitmap[2183] <= 1'b0;
		bitmap[2184] <= 1'b0;
		bitmap[2185] <= 1'b0;
		bitmap[2186] <= 1'b0;
		bitmap[2187] <= 1'b0;
		bitmap[2188] <= 1'b0;
		bitmap[2189] <= 1'b0;
		bitmap[2190] <= 1'b0;
		bitmap[2191] <= 1'b0;
		bitmap[2192] <= 1'b0;
		bitmap[2193] <= 1'b0;
		bitmap[2194] <= 1'b1;
		bitmap[2195] <= 1'b1;
		bitmap[2196] <= 1'b1;
		bitmap[2197] <= 1'b1;
		bitmap[2198] <= 1'b0;
		bitmap[2199] <= 1'b0;
		bitmap[2200] <= 1'b0;
		bitmap[2201] <= 1'b0;
		bitmap[2202] <= 1'b0;
		bitmap[2203] <= 1'b0;
		bitmap[2204] <= 1'b0;
		bitmap[2205] <= 1'b0;
		bitmap[2206] <= 1'b0;
		bitmap[2207] <= 1'b0;
		bitmap[2208] <= 1'b0;
		bitmap[2209] <= 1'b0;
		bitmap[2210] <= 1'b1;
		bitmap[2211] <= 1'b0;
		bitmap[2212] <= 1'b0;
		bitmap[2213] <= 1'b0;
		bitmap[2214] <= 1'b0;
		bitmap[2215] <= 1'b0;
		bitmap[2216] <= 1'b0;
		bitmap[2217] <= 1'b0;
		bitmap[2218] <= 1'b0;
		bitmap[2219] <= 1'b0;
		bitmap[2220] <= 1'b0;
		bitmap[2221] <= 1'b0;
		bitmap[2222] <= 1'b0;
		bitmap[2223] <= 1'b0;
		bitmap[2224] <= 1'b0;
		bitmap[2225] <= 1'b0;
		bitmap[2226] <= 1'b1;
		bitmap[2227] <= 1'b0;
		bitmap[2228] <= 1'b0;
		bitmap[2229] <= 1'b0;
		bitmap[2230] <= 1'b0;
		bitmap[2231] <= 1'b0;
		bitmap[2232] <= 1'b0;
		bitmap[2233] <= 1'b0;
		bitmap[2234] <= 1'b0;
		bitmap[2235] <= 1'b0;
		bitmap[2236] <= 1'b0;
		bitmap[2237] <= 1'b0;
		bitmap[2238] <= 1'b0;
		bitmap[2239] <= 1'b0;
		bitmap[2240] <= 1'b0;
		bitmap[2241] <= 1'b0;
		bitmap[2242] <= 1'b1;
		bitmap[2243] <= 1'b1;
		bitmap[2244] <= 1'b1;
		bitmap[2245] <= 1'b1;
		bitmap[2246] <= 1'b0;
		bitmap[2247] <= 1'b0;
		bitmap[2248] <= 1'b0;
		bitmap[2249] <= 1'b0;
		bitmap[2250] <= 1'b0;
		bitmap[2251] <= 1'b0;
		bitmap[2252] <= 1'b0;
		bitmap[2253] <= 1'b0;
		bitmap[2254] <= 1'b0;
		bitmap[2255] <= 1'b0;
		bitmap[2256] <= 1'b0;
		bitmap[2257] <= 1'b0;
		bitmap[2258] <= 1'b1;
		bitmap[2259] <= 1'b0;
		bitmap[2260] <= 1'b0;
		bitmap[2261] <= 1'b1;
		bitmap[2262] <= 1'b0;
		bitmap[2263] <= 1'b0;
		bitmap[2264] <= 1'b0;
		bitmap[2265] <= 1'b0;
		bitmap[2266] <= 1'b0;
		bitmap[2267] <= 1'b0;
		bitmap[2268] <= 1'b0;
		bitmap[2269] <= 1'b0;
		bitmap[2270] <= 1'b0;
		bitmap[2271] <= 1'b0;
		bitmap[2272] <= 1'b0;
		bitmap[2273] <= 1'b0;
		bitmap[2274] <= 1'b1;
		bitmap[2275] <= 1'b1;
		bitmap[2276] <= 1'b1;
		bitmap[2277] <= 1'b1;
		bitmap[2278] <= 1'b0;
		bitmap[2279] <= 1'b0;
		bitmap[2280] <= 1'b0;
		bitmap[2281] <= 1'b0;
		bitmap[2282] <= 1'b0;
		bitmap[2283] <= 1'b0;
		bitmap[2284] <= 1'b0;
		bitmap[2285] <= 1'b0;
		bitmap[2286] <= 1'b0;
		bitmap[2287] <= 1'b0;
		bitmap[2288] <= 1'b0;
		bitmap[2289] <= 1'b0;
		bitmap[2290] <= 1'b0;
		bitmap[2291] <= 1'b0;
		bitmap[2292] <= 1'b0;
		bitmap[2293] <= 1'b0;
		bitmap[2294] <= 1'b0;
		bitmap[2295] <= 1'b0;
		bitmap[2296] <= 1'b0;
		bitmap[2297] <= 1'b0;
		bitmap[2298] <= 1'b0;
		bitmap[2299] <= 1'b0;
		bitmap[2300] <= 1'b0;
		bitmap[2301] <= 1'b0;
		bitmap[2302] <= 1'b0;
		bitmap[2303] <= 1'b0;
		bitmap[2304] <= 1'b0;
		bitmap[2305] <= 1'b0;
		bitmap[2306] <= 1'b0;
		bitmap[2307] <= 1'b0;
		bitmap[2308] <= 1'b0;
		bitmap[2309] <= 1'b0;
		bitmap[2310] <= 1'b0;
		bitmap[2311] <= 1'b0;
		bitmap[2312] <= 1'b0;
		bitmap[2313] <= 1'b0;
		bitmap[2314] <= 1'b0;
		bitmap[2315] <= 1'b0;
		bitmap[2316] <= 1'b0;
		bitmap[2317] <= 1'b0;
		bitmap[2318] <= 1'b0;
		bitmap[2319] <= 1'b0;
		bitmap[2320] <= 1'b0;
		bitmap[2321] <= 1'b0;
		bitmap[2322] <= 1'b1;
		bitmap[2323] <= 1'b1;
		bitmap[2324] <= 1'b1;
		bitmap[2325] <= 1'b1;
		bitmap[2326] <= 1'b0;
		bitmap[2327] <= 1'b0;
		bitmap[2328] <= 1'b0;
		bitmap[2329] <= 1'b0;
		bitmap[2330] <= 1'b0;
		bitmap[2331] <= 1'b0;
		bitmap[2332] <= 1'b1;
		bitmap[2333] <= 1'b0;
		bitmap[2334] <= 1'b0;
		bitmap[2335] <= 1'b0;
		bitmap[2336] <= 1'b0;
		bitmap[2337] <= 1'b0;
		bitmap[2338] <= 1'b1;
		bitmap[2339] <= 1'b0;
		bitmap[2340] <= 1'b0;
		bitmap[2341] <= 1'b0;
		bitmap[2342] <= 1'b0;
		bitmap[2343] <= 1'b0;
		bitmap[2344] <= 1'b0;
		bitmap[2345] <= 1'b0;
		bitmap[2346] <= 1'b0;
		bitmap[2347] <= 1'b1;
		bitmap[2348] <= 1'b1;
		bitmap[2349] <= 1'b0;
		bitmap[2350] <= 1'b0;
		bitmap[2351] <= 1'b0;
		bitmap[2352] <= 1'b0;
		bitmap[2353] <= 1'b0;
		bitmap[2354] <= 1'b1;
		bitmap[2355] <= 1'b0;
		bitmap[2356] <= 1'b0;
		bitmap[2357] <= 1'b0;
		bitmap[2358] <= 1'b0;
		bitmap[2359] <= 1'b0;
		bitmap[2360] <= 1'b0;
		bitmap[2361] <= 1'b0;
		bitmap[2362] <= 1'b1;
		bitmap[2363] <= 1'b0;
		bitmap[2364] <= 1'b1;
		bitmap[2365] <= 1'b0;
		bitmap[2366] <= 1'b0;
		bitmap[2367] <= 1'b0;
		bitmap[2368] <= 1'b0;
		bitmap[2369] <= 1'b0;
		bitmap[2370] <= 1'b1;
		bitmap[2371] <= 1'b1;
		bitmap[2372] <= 1'b1;
		bitmap[2373] <= 1'b1;
		bitmap[2374] <= 1'b0;
		bitmap[2375] <= 1'b0;
		bitmap[2376] <= 1'b0;
		bitmap[2377] <= 1'b0;
		bitmap[2378] <= 1'b0;
		bitmap[2379] <= 1'b0;
		bitmap[2380] <= 1'b1;
		bitmap[2381] <= 1'b0;
		bitmap[2382] <= 1'b0;
		bitmap[2383] <= 1'b0;
		bitmap[2384] <= 1'b0;
		bitmap[2385] <= 1'b0;
		bitmap[2386] <= 1'b0;
		bitmap[2387] <= 1'b0;
		bitmap[2388] <= 1'b0;
		bitmap[2389] <= 1'b1;
		bitmap[2390] <= 1'b0;
		bitmap[2391] <= 1'b0;
		bitmap[2392] <= 1'b0;
		bitmap[2393] <= 1'b0;
		bitmap[2394] <= 1'b0;
		bitmap[2395] <= 1'b0;
		bitmap[2396] <= 1'b1;
		bitmap[2397] <= 1'b0;
		bitmap[2398] <= 1'b0;
		bitmap[2399] <= 1'b0;
		bitmap[2400] <= 1'b0;
		bitmap[2401] <= 1'b0;
		bitmap[2402] <= 1'b1;
		bitmap[2403] <= 1'b1;
		bitmap[2404] <= 1'b1;
		bitmap[2405] <= 1'b1;
		bitmap[2406] <= 1'b0;
		bitmap[2407] <= 1'b0;
		bitmap[2408] <= 1'b0;
		bitmap[2409] <= 1'b0;
		bitmap[2410] <= 1'b1;
		bitmap[2411] <= 1'b1;
		bitmap[2412] <= 1'b1;
		bitmap[2413] <= 1'b1;
		bitmap[2414] <= 1'b0;
		bitmap[2415] <= 1'b0;
		bitmap[2416] <= 1'b0;
		bitmap[2417] <= 1'b0;
		bitmap[2418] <= 1'b0;
		bitmap[2419] <= 1'b0;
		bitmap[2420] <= 1'b0;
		bitmap[2421] <= 1'b0;
		bitmap[2422] <= 1'b0;
		bitmap[2423] <= 1'b0;
		bitmap[2424] <= 1'b0;
		bitmap[2425] <= 1'b0;
		bitmap[2426] <= 1'b0;
		bitmap[2427] <= 1'b0;
		bitmap[2428] <= 1'b0;
		bitmap[2429] <= 1'b0;
		bitmap[2430] <= 1'b0;
		bitmap[2431] <= 1'b0;
		bitmap[2432] <= 1'b0;
		bitmap[2433] <= 1'b0;
		bitmap[2434] <= 1'b0;
		bitmap[2435] <= 1'b0;
		bitmap[2436] <= 1'b0;
		bitmap[2437] <= 1'b0;
		bitmap[2438] <= 1'b0;
		bitmap[2439] <= 1'b0;
		bitmap[2440] <= 1'b0;
		bitmap[2441] <= 1'b0;
		bitmap[2442] <= 1'b0;
		bitmap[2443] <= 1'b0;
		bitmap[2444] <= 1'b0;
		bitmap[2445] <= 1'b0;
		bitmap[2446] <= 1'b0;
		bitmap[2447] <= 1'b0;
		bitmap[2448] <= 1'b0;
		bitmap[2449] <= 1'b0;
		bitmap[2450] <= 1'b0;
		bitmap[2451] <= 1'b1;
		bitmap[2452] <= 1'b1;
		bitmap[2453] <= 1'b0;
		bitmap[2454] <= 1'b0;
		bitmap[2455] <= 1'b0;
		bitmap[2456] <= 1'b0;
		bitmap[2457] <= 1'b0;
		bitmap[2458] <= 1'b0;
		bitmap[2459] <= 1'b0;
		bitmap[2460] <= 1'b0;
		bitmap[2461] <= 1'b0;
		bitmap[2462] <= 1'b0;
		bitmap[2463] <= 1'b0;
		bitmap[2464] <= 1'b0;
		bitmap[2465] <= 1'b0;
		bitmap[2466] <= 1'b1;
		bitmap[2467] <= 1'b0;
		bitmap[2468] <= 1'b0;
		bitmap[2469] <= 1'b1;
		bitmap[2470] <= 1'b0;
		bitmap[2471] <= 1'b0;
		bitmap[2472] <= 1'b0;
		bitmap[2473] <= 1'b0;
		bitmap[2474] <= 1'b0;
		bitmap[2475] <= 1'b0;
		bitmap[2476] <= 1'b0;
		bitmap[2477] <= 1'b0;
		bitmap[2478] <= 1'b0;
		bitmap[2479] <= 1'b0;
		bitmap[2480] <= 1'b0;
		bitmap[2481] <= 1'b0;
		bitmap[2482] <= 1'b0;
		bitmap[2483] <= 1'b0;
		bitmap[2484] <= 1'b0;
		bitmap[2485] <= 1'b1;
		bitmap[2486] <= 1'b0;
		bitmap[2487] <= 1'b0;
		bitmap[2488] <= 1'b0;
		bitmap[2489] <= 1'b0;
		bitmap[2490] <= 1'b0;
		bitmap[2491] <= 1'b0;
		bitmap[2492] <= 1'b0;
		bitmap[2493] <= 1'b0;
		bitmap[2494] <= 1'b0;
		bitmap[2495] <= 1'b0;
		bitmap[2496] <= 1'b0;
		bitmap[2497] <= 1'b0;
		bitmap[2498] <= 1'b0;
		bitmap[2499] <= 1'b0;
		bitmap[2500] <= 1'b1;
		bitmap[2501] <= 1'b0;
		bitmap[2502] <= 1'b0;
		bitmap[2503] <= 1'b0;
		bitmap[2504] <= 1'b0;
		bitmap[2505] <= 1'b0;
		bitmap[2506] <= 1'b0;
		bitmap[2507] <= 1'b0;
		bitmap[2508] <= 1'b0;
		bitmap[2509] <= 1'b0;
		bitmap[2510] <= 1'b0;
		bitmap[2511] <= 1'b0;
		bitmap[2512] <= 1'b0;
		bitmap[2513] <= 1'b0;
		bitmap[2514] <= 1'b0;
		bitmap[2515] <= 1'b1;
		bitmap[2516] <= 1'b0;
		bitmap[2517] <= 1'b0;
		bitmap[2518] <= 1'b0;
		bitmap[2519] <= 1'b0;
		bitmap[2520] <= 1'b0;
		bitmap[2521] <= 1'b0;
		bitmap[2522] <= 1'b0;
		bitmap[2523] <= 1'b0;
		bitmap[2524] <= 1'b0;
		bitmap[2525] <= 1'b0;
		bitmap[2526] <= 1'b0;
		bitmap[2527] <= 1'b0;
		bitmap[2528] <= 1'b0;
		bitmap[2529] <= 1'b0;
		bitmap[2530] <= 1'b1;
		bitmap[2531] <= 1'b1;
		bitmap[2532] <= 1'b1;
		bitmap[2533] <= 1'b1;
		bitmap[2534] <= 1'b0;
		bitmap[2535] <= 1'b0;
		bitmap[2536] <= 1'b0;
		bitmap[2537] <= 1'b0;
		bitmap[2538] <= 1'b0;
		bitmap[2539] <= 1'b0;
		bitmap[2540] <= 1'b0;
		bitmap[2541] <= 1'b0;
		bitmap[2542] <= 1'b0;
		bitmap[2543] <= 1'b0;
		bitmap[2544] <= 1'b0;
		bitmap[2545] <= 1'b0;
		bitmap[2546] <= 1'b0;
		bitmap[2547] <= 1'b0;
		bitmap[2548] <= 1'b0;
		bitmap[2549] <= 1'b0;
		bitmap[2550] <= 1'b0;
		bitmap[2551] <= 1'b0;
		bitmap[2552] <= 1'b0;
		bitmap[2553] <= 1'b0;
		bitmap[2554] <= 1'b0;
		bitmap[2555] <= 1'b0;
		bitmap[2556] <= 1'b0;
		bitmap[2557] <= 1'b0;
		bitmap[2558] <= 1'b0;
		bitmap[2559] <= 1'b0;
		bitmap[2560] <= 1'b0;
		bitmap[2561] <= 1'b0;
		bitmap[2562] <= 1'b0;
		bitmap[2563] <= 1'b0;
		bitmap[2564] <= 1'b0;
		bitmap[2565] <= 1'b0;
		bitmap[2566] <= 1'b0;
		bitmap[2567] <= 1'b0;
		bitmap[2568] <= 1'b0;
		bitmap[2569] <= 1'b0;
		bitmap[2570] <= 1'b0;
		bitmap[2571] <= 1'b0;
		bitmap[2572] <= 1'b0;
		bitmap[2573] <= 1'b0;
		bitmap[2574] <= 1'b0;
		bitmap[2575] <= 1'b0;
		bitmap[2576] <= 1'b0;
		bitmap[2577] <= 1'b0;
		bitmap[2578] <= 1'b0;
		bitmap[2579] <= 1'b0;
		bitmap[2580] <= 1'b1;
		bitmap[2581] <= 1'b0;
		bitmap[2582] <= 1'b0;
		bitmap[2583] <= 1'b0;
		bitmap[2584] <= 1'b0;
		bitmap[2585] <= 1'b0;
		bitmap[2586] <= 1'b1;
		bitmap[2587] <= 1'b1;
		bitmap[2588] <= 1'b1;
		bitmap[2589] <= 1'b1;
		bitmap[2590] <= 1'b0;
		bitmap[2591] <= 1'b0;
		bitmap[2592] <= 1'b0;
		bitmap[2593] <= 1'b0;
		bitmap[2594] <= 1'b0;
		bitmap[2595] <= 1'b1;
		bitmap[2596] <= 1'b1;
		bitmap[2597] <= 1'b0;
		bitmap[2598] <= 1'b0;
		bitmap[2599] <= 1'b0;
		bitmap[2600] <= 1'b0;
		bitmap[2601] <= 1'b0;
		bitmap[2602] <= 1'b1;
		bitmap[2603] <= 1'b0;
		bitmap[2604] <= 1'b0;
		bitmap[2605] <= 1'b1;
		bitmap[2606] <= 1'b0;
		bitmap[2607] <= 1'b0;
		bitmap[2608] <= 1'b0;
		bitmap[2609] <= 1'b0;
		bitmap[2610] <= 1'b1;
		bitmap[2611] <= 1'b0;
		bitmap[2612] <= 1'b1;
		bitmap[2613] <= 1'b0;
		bitmap[2614] <= 1'b0;
		bitmap[2615] <= 1'b0;
		bitmap[2616] <= 1'b0;
		bitmap[2617] <= 1'b0;
		bitmap[2618] <= 1'b1;
		bitmap[2619] <= 1'b0;
		bitmap[2620] <= 1'b0;
		bitmap[2621] <= 1'b1;
		bitmap[2622] <= 1'b0;
		bitmap[2623] <= 1'b0;
		bitmap[2624] <= 1'b0;
		bitmap[2625] <= 1'b0;
		bitmap[2626] <= 1'b0;
		bitmap[2627] <= 1'b0;
		bitmap[2628] <= 1'b1;
		bitmap[2629] <= 1'b0;
		bitmap[2630] <= 1'b0;
		bitmap[2631] <= 1'b0;
		bitmap[2632] <= 1'b0;
		bitmap[2633] <= 1'b0;
		bitmap[2634] <= 1'b1;
		bitmap[2635] <= 1'b0;
		bitmap[2636] <= 1'b0;
		bitmap[2637] <= 1'b1;
		bitmap[2638] <= 1'b0;
		bitmap[2639] <= 1'b0;
		bitmap[2640] <= 1'b0;
		bitmap[2641] <= 1'b0;
		bitmap[2642] <= 1'b0;
		bitmap[2643] <= 1'b0;
		bitmap[2644] <= 1'b1;
		bitmap[2645] <= 1'b0;
		bitmap[2646] <= 1'b0;
		bitmap[2647] <= 1'b0;
		bitmap[2648] <= 1'b0;
		bitmap[2649] <= 1'b0;
		bitmap[2650] <= 1'b1;
		bitmap[2651] <= 1'b0;
		bitmap[2652] <= 1'b0;
		bitmap[2653] <= 1'b1;
		bitmap[2654] <= 1'b0;
		bitmap[2655] <= 1'b0;
		bitmap[2656] <= 1'b0;
		bitmap[2657] <= 1'b0;
		bitmap[2658] <= 1'b1;
		bitmap[2659] <= 1'b1;
		bitmap[2660] <= 1'b1;
		bitmap[2661] <= 1'b1;
		bitmap[2662] <= 1'b0;
		bitmap[2663] <= 1'b0;
		bitmap[2664] <= 1'b0;
		bitmap[2665] <= 1'b0;
		bitmap[2666] <= 1'b1;
		bitmap[2667] <= 1'b1;
		bitmap[2668] <= 1'b1;
		bitmap[2669] <= 1'b1;
		bitmap[2670] <= 1'b0;
		bitmap[2671] <= 1'b0;
		bitmap[2672] <= 1'b0;
		bitmap[2673] <= 1'b0;
		bitmap[2674] <= 1'b0;
		bitmap[2675] <= 1'b0;
		bitmap[2676] <= 1'b0;
		bitmap[2677] <= 1'b0;
		bitmap[2678] <= 1'b0;
		bitmap[2679] <= 1'b0;
		bitmap[2680] <= 1'b0;
		bitmap[2681] <= 1'b0;
		bitmap[2682] <= 1'b0;
		bitmap[2683] <= 1'b0;
		bitmap[2684] <= 1'b0;
		bitmap[2685] <= 1'b0;
		bitmap[2686] <= 1'b0;
		bitmap[2687] <= 1'b0;
		bitmap[2688] <= 1'b0;
		bitmap[2689] <= 1'b0;
		bitmap[2690] <= 1'b0;
		bitmap[2691] <= 1'b0;
		bitmap[2692] <= 1'b0;
		bitmap[2693] <= 1'b0;
		bitmap[2694] <= 1'b0;
		bitmap[2695] <= 1'b0;
		bitmap[2696] <= 1'b0;
		bitmap[2697] <= 1'b0;
		bitmap[2698] <= 1'b0;
		bitmap[2699] <= 1'b0;
		bitmap[2700] <= 1'b0;
		bitmap[2701] <= 1'b0;
		bitmap[2702] <= 1'b0;
		bitmap[2703] <= 1'b0;
		bitmap[2704] <= 1'b0;
		bitmap[2705] <= 1'b0;
		bitmap[2706] <= 1'b0;
		bitmap[2707] <= 1'b1;
		bitmap[2708] <= 1'b1;
		bitmap[2709] <= 1'b0;
		bitmap[2710] <= 1'b0;
		bitmap[2711] <= 1'b0;
		bitmap[2712] <= 1'b0;
		bitmap[2713] <= 1'b0;
		bitmap[2714] <= 1'b0;
		bitmap[2715] <= 1'b0;
		bitmap[2716] <= 1'b1;
		bitmap[2717] <= 1'b1;
		bitmap[2718] <= 1'b0;
		bitmap[2719] <= 1'b0;
		bitmap[2720] <= 1'b0;
		bitmap[2721] <= 1'b0;
		bitmap[2722] <= 1'b1;
		bitmap[2723] <= 1'b0;
		bitmap[2724] <= 1'b0;
		bitmap[2725] <= 1'b1;
		bitmap[2726] <= 1'b0;
		bitmap[2727] <= 1'b0;
		bitmap[2728] <= 1'b0;
		bitmap[2729] <= 1'b0;
		bitmap[2730] <= 1'b0;
		bitmap[2731] <= 1'b1;
		bitmap[2732] <= 1'b0;
		bitmap[2733] <= 1'b1;
		bitmap[2734] <= 1'b0;
		bitmap[2735] <= 1'b0;
		bitmap[2736] <= 1'b0;
		bitmap[2737] <= 1'b0;
		bitmap[2738] <= 1'b0;
		bitmap[2739] <= 1'b0;
		bitmap[2740] <= 1'b0;
		bitmap[2741] <= 1'b1;
		bitmap[2742] <= 1'b0;
		bitmap[2743] <= 1'b0;
		bitmap[2744] <= 1'b0;
		bitmap[2745] <= 1'b0;
		bitmap[2746] <= 1'b1;
		bitmap[2747] <= 1'b0;
		bitmap[2748] <= 1'b0;
		bitmap[2749] <= 1'b1;
		bitmap[2750] <= 1'b0;
		bitmap[2751] <= 1'b0;
		bitmap[2752] <= 1'b0;
		bitmap[2753] <= 1'b0;
		bitmap[2754] <= 1'b0;
		bitmap[2755] <= 1'b0;
		bitmap[2756] <= 1'b1;
		bitmap[2757] <= 1'b0;
		bitmap[2758] <= 1'b0;
		bitmap[2759] <= 1'b0;
		bitmap[2760] <= 1'b0;
		bitmap[2761] <= 1'b0;
		bitmap[2762] <= 1'b1;
		bitmap[2763] <= 1'b1;
		bitmap[2764] <= 1'b1;
		bitmap[2765] <= 1'b1;
		bitmap[2766] <= 1'b1;
		bitmap[2767] <= 1'b0;
		bitmap[2768] <= 1'b0;
		bitmap[2769] <= 1'b0;
		bitmap[2770] <= 1'b0;
		bitmap[2771] <= 1'b1;
		bitmap[2772] <= 1'b0;
		bitmap[2773] <= 1'b0;
		bitmap[2774] <= 1'b0;
		bitmap[2775] <= 1'b0;
		bitmap[2776] <= 1'b0;
		bitmap[2777] <= 1'b0;
		bitmap[2778] <= 1'b0;
		bitmap[2779] <= 1'b0;
		bitmap[2780] <= 1'b0;
		bitmap[2781] <= 1'b1;
		bitmap[2782] <= 1'b0;
		bitmap[2783] <= 1'b0;
		bitmap[2784] <= 1'b0;
		bitmap[2785] <= 1'b0;
		bitmap[2786] <= 1'b1;
		bitmap[2787] <= 1'b1;
		bitmap[2788] <= 1'b1;
		bitmap[2789] <= 1'b1;
		bitmap[2790] <= 1'b0;
		bitmap[2791] <= 1'b0;
		bitmap[2792] <= 1'b0;
		bitmap[2793] <= 1'b0;
		bitmap[2794] <= 1'b0;
		bitmap[2795] <= 1'b0;
		bitmap[2796] <= 1'b0;
		bitmap[2797] <= 1'b1;
		bitmap[2798] <= 1'b0;
		bitmap[2799] <= 1'b0;
		bitmap[2800] <= 1'b0;
		bitmap[2801] <= 1'b0;
		bitmap[2802] <= 1'b0;
		bitmap[2803] <= 1'b0;
		bitmap[2804] <= 1'b0;
		bitmap[2805] <= 1'b0;
		bitmap[2806] <= 1'b0;
		bitmap[2807] <= 1'b0;
		bitmap[2808] <= 1'b0;
		bitmap[2809] <= 1'b0;
		bitmap[2810] <= 1'b0;
		bitmap[2811] <= 1'b0;
		bitmap[2812] <= 1'b0;
		bitmap[2813] <= 1'b0;
		bitmap[2814] <= 1'b0;
		bitmap[2815] <= 1'b0;
		bitmap[2816] <= 1'b0;
		bitmap[2817] <= 1'b0;
		bitmap[2818] <= 1'b0;
		bitmap[2819] <= 1'b0;
		bitmap[2820] <= 1'b0;
		bitmap[2821] <= 1'b0;
		bitmap[2822] <= 1'b0;
		bitmap[2823] <= 1'b0;
		bitmap[2824] <= 1'b0;
		bitmap[2825] <= 1'b0;
		bitmap[2826] <= 1'b0;
		bitmap[2827] <= 1'b0;
		bitmap[2828] <= 1'b0;
		bitmap[2829] <= 1'b0;
		bitmap[2830] <= 1'b0;
		bitmap[2831] <= 1'b0;
		bitmap[2832] <= 1'b0;
		bitmap[2833] <= 1'b0;
		bitmap[2834] <= 1'b0;
		bitmap[2835] <= 1'b1;
		bitmap[2836] <= 1'b1;
		bitmap[2837] <= 1'b0;
		bitmap[2838] <= 1'b0;
		bitmap[2839] <= 1'b0;
		bitmap[2840] <= 1'b0;
		bitmap[2841] <= 1'b0;
		bitmap[2842] <= 1'b1;
		bitmap[2843] <= 1'b1;
		bitmap[2844] <= 1'b1;
		bitmap[2845] <= 1'b1;
		bitmap[2846] <= 1'b0;
		bitmap[2847] <= 1'b0;
		bitmap[2848] <= 1'b0;
		bitmap[2849] <= 1'b0;
		bitmap[2850] <= 1'b1;
		bitmap[2851] <= 1'b0;
		bitmap[2852] <= 1'b0;
		bitmap[2853] <= 1'b1;
		bitmap[2854] <= 1'b0;
		bitmap[2855] <= 1'b0;
		bitmap[2856] <= 1'b0;
		bitmap[2857] <= 1'b0;
		bitmap[2858] <= 1'b1;
		bitmap[2859] <= 1'b0;
		bitmap[2860] <= 1'b0;
		bitmap[2861] <= 1'b1;
		bitmap[2862] <= 1'b0;
		bitmap[2863] <= 1'b0;
		bitmap[2864] <= 1'b0;
		bitmap[2865] <= 1'b0;
		bitmap[2866] <= 1'b0;
		bitmap[2867] <= 1'b0;
		bitmap[2868] <= 1'b0;
		bitmap[2869] <= 1'b1;
		bitmap[2870] <= 1'b0;
		bitmap[2871] <= 1'b0;
		bitmap[2872] <= 1'b0;
		bitmap[2873] <= 1'b0;
		bitmap[2874] <= 1'b1;
		bitmap[2875] <= 1'b0;
		bitmap[2876] <= 1'b0;
		bitmap[2877] <= 1'b1;
		bitmap[2878] <= 1'b0;
		bitmap[2879] <= 1'b0;
		bitmap[2880] <= 1'b0;
		bitmap[2881] <= 1'b0;
		bitmap[2882] <= 1'b0;
		bitmap[2883] <= 1'b0;
		bitmap[2884] <= 1'b1;
		bitmap[2885] <= 1'b0;
		bitmap[2886] <= 1'b0;
		bitmap[2887] <= 1'b0;
		bitmap[2888] <= 1'b0;
		bitmap[2889] <= 1'b0;
		bitmap[2890] <= 1'b1;
		bitmap[2891] <= 1'b0;
		bitmap[2892] <= 1'b0;
		bitmap[2893] <= 1'b1;
		bitmap[2894] <= 1'b0;
		bitmap[2895] <= 1'b0;
		bitmap[2896] <= 1'b0;
		bitmap[2897] <= 1'b0;
		bitmap[2898] <= 1'b0;
		bitmap[2899] <= 1'b1;
		bitmap[2900] <= 1'b0;
		bitmap[2901] <= 1'b0;
		bitmap[2902] <= 1'b0;
		bitmap[2903] <= 1'b0;
		bitmap[2904] <= 1'b0;
		bitmap[2905] <= 1'b0;
		bitmap[2906] <= 1'b1;
		bitmap[2907] <= 1'b0;
		bitmap[2908] <= 1'b0;
		bitmap[2909] <= 1'b1;
		bitmap[2910] <= 1'b0;
		bitmap[2911] <= 1'b0;
		bitmap[2912] <= 1'b0;
		bitmap[2913] <= 1'b0;
		bitmap[2914] <= 1'b1;
		bitmap[2915] <= 1'b1;
		bitmap[2916] <= 1'b1;
		bitmap[2917] <= 1'b1;
		bitmap[2918] <= 1'b0;
		bitmap[2919] <= 1'b0;
		bitmap[2920] <= 1'b0;
		bitmap[2921] <= 1'b0;
		bitmap[2922] <= 1'b1;
		bitmap[2923] <= 1'b1;
		bitmap[2924] <= 1'b1;
		bitmap[2925] <= 1'b1;
		bitmap[2926] <= 1'b0;
		bitmap[2927] <= 1'b0;
		bitmap[2928] <= 1'b0;
		bitmap[2929] <= 1'b0;
		bitmap[2930] <= 1'b0;
		bitmap[2931] <= 1'b0;
		bitmap[2932] <= 1'b0;
		bitmap[2933] <= 1'b0;
		bitmap[2934] <= 1'b0;
		bitmap[2935] <= 1'b0;
		bitmap[2936] <= 1'b0;
		bitmap[2937] <= 1'b0;
		bitmap[2938] <= 1'b0;
		bitmap[2939] <= 1'b0;
		bitmap[2940] <= 1'b0;
		bitmap[2941] <= 1'b0;
		bitmap[2942] <= 1'b0;
		bitmap[2943] <= 1'b0;
		bitmap[2944] <= 1'b0;
		bitmap[2945] <= 1'b0;
		bitmap[2946] <= 1'b0;
		bitmap[2947] <= 1'b0;
		bitmap[2948] <= 1'b0;
		bitmap[2949] <= 1'b0;
		bitmap[2950] <= 1'b0;
		bitmap[2951] <= 1'b0;
		bitmap[2952] <= 1'b0;
		bitmap[2953] <= 1'b0;
		bitmap[2954] <= 1'b0;
		bitmap[2955] <= 1'b0;
		bitmap[2956] <= 1'b0;
		bitmap[2957] <= 1'b0;
		bitmap[2958] <= 1'b0;
		bitmap[2959] <= 1'b0;
		bitmap[2960] <= 1'b0;
		bitmap[2961] <= 1'b0;
		bitmap[2962] <= 1'b0;
		bitmap[2963] <= 1'b0;
		bitmap[2964] <= 1'b1;
		bitmap[2965] <= 1'b1;
		bitmap[2966] <= 1'b0;
		bitmap[2967] <= 1'b0;
		bitmap[2968] <= 1'b0;
		bitmap[2969] <= 1'b0;
		bitmap[2970] <= 1'b1;
		bitmap[2971] <= 1'b1;
		bitmap[2972] <= 1'b1;
		bitmap[2973] <= 1'b1;
		bitmap[2974] <= 1'b0;
		bitmap[2975] <= 1'b0;
		bitmap[2976] <= 1'b0;
		bitmap[2977] <= 1'b0;
		bitmap[2978] <= 1'b0;
		bitmap[2979] <= 1'b1;
		bitmap[2980] <= 1'b0;
		bitmap[2981] <= 1'b1;
		bitmap[2982] <= 1'b0;
		bitmap[2983] <= 1'b0;
		bitmap[2984] <= 1'b0;
		bitmap[2985] <= 1'b0;
		bitmap[2986] <= 1'b1;
		bitmap[2987] <= 1'b0;
		bitmap[2988] <= 1'b0;
		bitmap[2989] <= 1'b1;
		bitmap[2990] <= 1'b0;
		bitmap[2991] <= 1'b0;
		bitmap[2992] <= 1'b0;
		bitmap[2993] <= 1'b0;
		bitmap[2994] <= 1'b1;
		bitmap[2995] <= 1'b0;
		bitmap[2996] <= 1'b0;
		bitmap[2997] <= 1'b1;
		bitmap[2998] <= 1'b0;
		bitmap[2999] <= 1'b0;
		bitmap[3000] <= 1'b0;
		bitmap[3001] <= 1'b0;
		bitmap[3002] <= 1'b1;
		bitmap[3003] <= 1'b0;
		bitmap[3004] <= 1'b0;
		bitmap[3005] <= 1'b1;
		bitmap[3006] <= 1'b0;
		bitmap[3007] <= 1'b0;
		bitmap[3008] <= 1'b0;
		bitmap[3009] <= 1'b0;
		bitmap[3010] <= 1'b1;
		bitmap[3011] <= 1'b1;
		bitmap[3012] <= 1'b1;
		bitmap[3013] <= 1'b1;
		bitmap[3014] <= 1'b1;
		bitmap[3015] <= 1'b0;
		bitmap[3016] <= 1'b0;
		bitmap[3017] <= 1'b0;
		bitmap[3018] <= 1'b1;
		bitmap[3019] <= 1'b1;
		bitmap[3020] <= 1'b1;
		bitmap[3021] <= 1'b1;
		bitmap[3022] <= 1'b0;
		bitmap[3023] <= 1'b0;
		bitmap[3024] <= 1'b0;
		bitmap[3025] <= 1'b0;
		bitmap[3026] <= 1'b0;
		bitmap[3027] <= 1'b0;
		bitmap[3028] <= 1'b0;
		bitmap[3029] <= 1'b1;
		bitmap[3030] <= 1'b0;
		bitmap[3031] <= 1'b0;
		bitmap[3032] <= 1'b0;
		bitmap[3033] <= 1'b0;
		bitmap[3034] <= 1'b1;
		bitmap[3035] <= 1'b0;
		bitmap[3036] <= 1'b0;
		bitmap[3037] <= 1'b1;
		bitmap[3038] <= 1'b0;
		bitmap[3039] <= 1'b0;
		bitmap[3040] <= 1'b0;
		bitmap[3041] <= 1'b0;
		bitmap[3042] <= 1'b0;
		bitmap[3043] <= 1'b0;
		bitmap[3044] <= 1'b0;
		bitmap[3045] <= 1'b1;
		bitmap[3046] <= 1'b0;
		bitmap[3047] <= 1'b0;
		bitmap[3048] <= 1'b0;
		bitmap[3049] <= 1'b0;
		bitmap[3050] <= 1'b1;
		bitmap[3051] <= 1'b1;
		bitmap[3052] <= 1'b1;
		bitmap[3053] <= 1'b1;
		bitmap[3054] <= 1'b0;
		bitmap[3055] <= 1'b0;
		bitmap[3056] <= 1'b0;
		bitmap[3057] <= 1'b0;
		bitmap[3058] <= 1'b0;
		bitmap[3059] <= 1'b0;
		bitmap[3060] <= 1'b0;
		bitmap[3061] <= 1'b0;
		bitmap[3062] <= 1'b0;
		bitmap[3063] <= 1'b0;
		bitmap[3064] <= 1'b0;
		bitmap[3065] <= 1'b0;
		bitmap[3066] <= 1'b0;
		bitmap[3067] <= 1'b0;
		bitmap[3068] <= 1'b0;
		bitmap[3069] <= 1'b0;
		bitmap[3070] <= 1'b0;
		bitmap[3071] <= 1'b0;

		palette[0]  <= 12'b1111_1111_1111;
		palette[1]  <= 12'b0000_0000_0000;
		palette[2]  <= 12'b1111_0000_0000;
		palette[3]  <= 12'b0000_0000_0000;
		palette[4]  <= 12'b1111_1000_0000;
		palette[5]  <= 12'b0000_0000_0000;
		palette[6]  <= 12'b1111_1111_0000;
		palette[7]  <= 12'b0000_0000_0000;
		palette[8]  <= 12'b1000_1111_0000;
		palette[9]  <= 12'b0000_0000_0000;
		palette[10] <= 12'b0000_1111_0000;
		palette[11] <= 12'b0000_0000_0000;
		palette[12] <= 12'b0000_1111_1000;
		palette[13] <= 12'b0000_0000_0000;
		palette[14] <= 12'b0000_1111_1111;
		palette[15] <= 12'b0000_0000_0000;
		palette[16] <= 12'b0000_1000_1111;
		palette[17] <= 12'b0000_0000_0000;
		palette[18] <= 12'b0000_0000_1111;
		palette[19] <= 12'b0000_0000_0000;
		palette[20] <= 12'b1000_0000_1111;
		palette[21] <= 12'b0000_0000_0000;
		palette[22] <= 12'b1111_0000_1111;
		palette[23] <= 12'b0000_0000_0000;
	end

endmodule
