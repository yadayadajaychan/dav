module vga_top (
	input clk, // 50 MHz
	input rst,

	output logic hsync,
	output logic vsync,
	output logic [3:0] red,
	output logic [3:0] green,
	output logic [3:0] blue
);

	wire vgaclk;
	clock_divider divider1(clk, rst, vgaclk);
	reg [7:0] color;

	localparam BLK = 8'h00;
	localparam WHT = 8'hff;
	localparam RED = 8'he0;
	localparam BLU = 8'h03;
	reg [7:0] test_sprite [0:767];

	wire [9:0] hc_out;
	wire [9:0] vc_out;
	vga vga1(vgaclk, rst, color[7:5], color[4:2], color[1:0],
		hc_out, vc_out, hsync, vsync, red, green, blue);

	reg [9:0] i;
	always @(posedge vgaclk) begin
		color <= test_sprite[i];

		if (!rst || i >= 768) begin
			i <= 0;
		end else begin
			if (hc_out < 32) begin
				i <= i + 1;
			end
		end
	end

	always @(negedge rst) begin
		test_sprite[0] = BLK;
		test_sprite[1] = BLK;
		test_sprite[2] = BLK;
		test_sprite[3] = BLK;
		test_sprite[4] = BLK;
		test_sprite[5] = BLK;
		test_sprite[6] = BLK;
		test_sprite[7] = BLK;
		test_sprite[8] = BLK;
		test_sprite[9] = BLK;
		test_sprite[10] = BLK;
		test_sprite[11] = BLK;
		test_sprite[12] = BLK;
		test_sprite[13] = BLK;
		test_sprite[14] = BLK;
		test_sprite[15] = BLK;
		test_sprite[16] = BLK;
		test_sprite[17] = BLK;
		test_sprite[18] = BLK;
		test_sprite[19] = BLK;
		test_sprite[20] = BLK;
		test_sprite[21] = BLK;
		test_sprite[22] = BLK;
		test_sprite[23] = BLK;
		test_sprite[24] = BLK;
		test_sprite[25] = BLK;
		test_sprite[26] = BLK;
		test_sprite[27] = BLK;
		test_sprite[28] = BLK;
		test_sprite[29] = BLK;
		test_sprite[30] = BLK;
		test_sprite[31] = BLK;
		test_sprite[32] = BLK;
		test_sprite[33] = BLK;
		test_sprite[34] = BLK;
		test_sprite[35] = BLK;
		test_sprite[36] = BLK;
		test_sprite[37] = BLK;
		test_sprite[38] = BLK;
		test_sprite[39] = BLK;
		test_sprite[40] = BLK;
		test_sprite[41] = BLK;
		test_sprite[42] = BLK;
		test_sprite[43] = BLK;
		test_sprite[44] = BLK;
		test_sprite[45] = BLK;
		test_sprite[46] = BLK;
		test_sprite[47] = BLK;
		test_sprite[48] = BLK;
		test_sprite[49] = BLK;
		test_sprite[50] = BLK;
		test_sprite[51] = BLK;
		test_sprite[52] = BLK;
		test_sprite[53] = BLK;
		test_sprite[54] = BLK;
		test_sprite[55] = BLK;
		test_sprite[56] = BLK;
		test_sprite[57] = BLK;
		test_sprite[58] = BLK;
		test_sprite[59] = BLK;
		test_sprite[60] = BLK;
		test_sprite[61] = BLK;
		test_sprite[62] = BLK;
		test_sprite[63] = BLK;
		test_sprite[64] = BLK;
		test_sprite[65] = BLK;
		test_sprite[66] = BLK;
		test_sprite[67] = BLK;
		test_sprite[68] = BLK;
		test_sprite[69] = BLK;
		test_sprite[70] = BLK;
		test_sprite[71] = BLK;
		test_sprite[72] = BLK;
		test_sprite[73] = BLK;
		test_sprite[74] = BLK;
		test_sprite[75] = BLK;
		test_sprite[76] = BLK;
		test_sprite[77] = BLK;
		test_sprite[78] = BLK;
		test_sprite[79] = BLK;
		test_sprite[80] = BLK;
		test_sprite[81] = BLK;
		test_sprite[82] = BLK;
		test_sprite[83] = BLK;
		test_sprite[84] = BLK;
		test_sprite[85] = BLK;
		test_sprite[86] = BLK;
		test_sprite[87] = BLK;
		test_sprite[88] = BLK;
		test_sprite[89] = BLK;
		test_sprite[90] = BLK;
		test_sprite[91] = BLK;
		test_sprite[92] = BLK;
		test_sprite[93] = BLK;
		test_sprite[94] = BLK;
		test_sprite[95] = BLK;
		test_sprite[96] = BLK;
		test_sprite[97] = BLK;
		test_sprite[98] = BLK;
		test_sprite[99] = BLK;
		test_sprite[100] = BLK;
		test_sprite[101] = BLK;
		test_sprite[102] = BLK;
		test_sprite[103] = BLK;
		test_sprite[104] = BLK;
		test_sprite[105] = BLK;
		test_sprite[106] = BLK;
		test_sprite[107] = BLK;
		test_sprite[108] = BLK;
		test_sprite[109] = BLK;
		test_sprite[110] = BLK;
		test_sprite[111] = BLK;
		test_sprite[112] = BLK;
		test_sprite[113] = BLK;
		test_sprite[114] = BLK;
		test_sprite[115] = BLK;
		test_sprite[116] = BLK;
		test_sprite[117] = BLK;
		test_sprite[118] = BLK;
		test_sprite[119] = BLK;
		test_sprite[120] = BLK;
		test_sprite[121] = BLK;
		test_sprite[122] = BLK;
		test_sprite[123] = BLK;
		test_sprite[124] = BLK;
		test_sprite[125] = BLK;
		test_sprite[126] = BLK;
		test_sprite[127] = BLK;
		test_sprite[128] = BLK;
		test_sprite[129] = BLK;
		test_sprite[130] = BLK;
		test_sprite[131] = BLK;
		test_sprite[132] = BLK;
		test_sprite[133] = BLK;
		test_sprite[134] = BLK;
		test_sprite[135] = BLK;
		test_sprite[136] = BLK;
		test_sprite[137] = BLK;
		test_sprite[138] = BLK;
		test_sprite[139] = BLK;
		test_sprite[140] = BLK;
		test_sprite[141] = BLK;
		test_sprite[142] = BLK;
		test_sprite[143] = BLK;
		test_sprite[144] = BLK;
		test_sprite[145] = BLK;
		test_sprite[146] = BLK;
		test_sprite[147] = BLK;
		test_sprite[148] = BLK;
		test_sprite[149] = BLK;
		test_sprite[150] = BLK;
		test_sprite[151] = BLK;
		test_sprite[152] = BLK;
		test_sprite[153] = BLK;
		test_sprite[154] = BLK;
		test_sprite[155] = BLK;
		test_sprite[156] = BLK;
		test_sprite[157] = BLK;
		test_sprite[158] = BLK;
		test_sprite[159] = BLK;
		test_sprite[160] = BLK;
		test_sprite[161] = BLK;
		test_sprite[162] = BLK;
		test_sprite[163] = BLK;
		test_sprite[164] = BLK;
		test_sprite[165] = BLK;
		test_sprite[166] = BLK;
		test_sprite[167] = BLK;
		test_sprite[168] = BLK;
		test_sprite[169] = BLK;
		test_sprite[170] = BLK;
		test_sprite[171] = BLK;
		test_sprite[172] = BLK;
		test_sprite[173] = BLK;
		test_sprite[174] = RED;
		test_sprite[175] = RED;
		test_sprite[176] = RED;
		test_sprite[177] = RED;
		test_sprite[178] = BLK;
		test_sprite[179] = BLK;
		test_sprite[180] = BLK;
		test_sprite[181] = BLK;
		test_sprite[182] = BLK;
		test_sprite[183] = BLK;
		test_sprite[184] = BLK;
		test_sprite[185] = BLK;
		test_sprite[186] = BLK;
		test_sprite[187] = BLK;
		test_sprite[188] = BLK;
		test_sprite[189] = BLK;
		test_sprite[190] = BLK;
		test_sprite[191] = BLK;
		test_sprite[192] = BLK;
		test_sprite[193] = BLK;
		test_sprite[194] = BLK;
		test_sprite[195] = BLK;
		test_sprite[196] = BLK;
		test_sprite[197] = BLK;
		test_sprite[198] = BLK;
		test_sprite[199] = BLK;
		test_sprite[200] = BLK;
		test_sprite[201] = BLK;
		test_sprite[202] = BLK;
		test_sprite[203] = BLK;
		test_sprite[204] = RED;
		test_sprite[205] = RED;
		test_sprite[206] = RED;
		test_sprite[207] = RED;
		test_sprite[208] = RED;
		test_sprite[209] = RED;
		test_sprite[210] = RED;
		test_sprite[211] = RED;
		test_sprite[212] = BLK;
		test_sprite[213] = BLK;
		test_sprite[214] = BLK;
		test_sprite[215] = BLK;
		test_sprite[216] = BLK;
		test_sprite[217] = BLK;
		test_sprite[218] = BLK;
		test_sprite[219] = BLK;
		test_sprite[220] = BLK;
		test_sprite[221] = BLK;
		test_sprite[222] = BLK;
		test_sprite[223] = BLK;
		test_sprite[224] = BLK;
		test_sprite[225] = BLK;
		test_sprite[226] = BLK;
		test_sprite[227] = BLK;
		test_sprite[228] = BLK;
		test_sprite[229] = BLK;
		test_sprite[230] = BLK;
		test_sprite[231] = BLK;
		test_sprite[232] = BLK;
		test_sprite[233] = BLK;
		test_sprite[234] = BLK;
		test_sprite[235] = RED;
		test_sprite[236] = RED;
		test_sprite[237] = RED;
		test_sprite[238] = RED;
		test_sprite[239] = RED;
		test_sprite[240] = RED;
		test_sprite[241] = RED;
		test_sprite[242] = RED;
		test_sprite[243] = RED;
		test_sprite[244] = RED;
		test_sprite[245] = BLK;
		test_sprite[246] = BLK;
		test_sprite[247] = BLK;
		test_sprite[248] = BLK;
		test_sprite[249] = BLK;
		test_sprite[250] = BLK;
		test_sprite[251] = BLK;
		test_sprite[252] = BLK;
		test_sprite[253] = BLK;
		test_sprite[254] = BLK;
		test_sprite[255] = BLK;
		test_sprite[256] = BLK;
		test_sprite[257] = BLK;
		test_sprite[258] = BLK;
		test_sprite[259] = BLK;
		test_sprite[260] = BLK;
		test_sprite[261] = BLK;
		test_sprite[262] = BLK;
		test_sprite[263] = BLK;
		test_sprite[264] = BLK;
		test_sprite[265] = BLK;
		test_sprite[266] = RED;
		test_sprite[267] = RED;
		test_sprite[268] = RED;
		test_sprite[269] = WHT;
		test_sprite[270] = WHT;
		test_sprite[271] = RED;
		test_sprite[272] = RED;
		test_sprite[273] = RED;
		test_sprite[274] = RED;
		test_sprite[275] = WHT;
		test_sprite[276] = WHT;
		test_sprite[277] = RED;
		test_sprite[278] = BLK;
		test_sprite[279] = BLK;
		test_sprite[280] = BLK;
		test_sprite[281] = BLK;
		test_sprite[282] = BLK;
		test_sprite[283] = BLK;
		test_sprite[284] = BLK;
		test_sprite[285] = BLK;
		test_sprite[286] = BLK;
		test_sprite[287] = BLK;
		test_sprite[288] = BLK;
		test_sprite[289] = BLK;
		test_sprite[290] = BLK;
		test_sprite[291] = BLK;
		test_sprite[292] = BLK;
		test_sprite[293] = BLK;
		test_sprite[294] = BLK;
		test_sprite[295] = BLK;
		test_sprite[296] = BLK;
		test_sprite[297] = BLK;
		test_sprite[298] = RED;
		test_sprite[299] = RED;
		test_sprite[300] = WHT;
		test_sprite[301] = WHT;
		test_sprite[302] = WHT;
		test_sprite[303] = WHT;
		test_sprite[304] = RED;
		test_sprite[305] = RED;
		test_sprite[306] = WHT;
		test_sprite[307] = WHT;
		test_sprite[308] = WHT;
		test_sprite[309] = WHT;
		test_sprite[310] = BLK;
		test_sprite[311] = BLK;
		test_sprite[312] = BLK;
		test_sprite[313] = BLK;
		test_sprite[314] = BLK;
		test_sprite[315] = BLK;
		test_sprite[316] = BLK;
		test_sprite[317] = BLK;
		test_sprite[318] = BLK;
		test_sprite[319] = BLK;
		test_sprite[320] = BLK;
		test_sprite[321] = BLK;
		test_sprite[322] = BLK;
		test_sprite[323] = BLK;
		test_sprite[324] = BLK;
		test_sprite[325] = BLK;
		test_sprite[326] = BLK;
		test_sprite[327] = BLK;
		test_sprite[328] = BLK;
		test_sprite[329] = BLK;
		test_sprite[330] = RED;
		test_sprite[331] = RED;
		test_sprite[332] = WHT;
		test_sprite[333] = WHT;
		test_sprite[334] = BLU;
		test_sprite[335] = BLU;
		test_sprite[336] = RED;
		test_sprite[337] = RED;
		test_sprite[338] = WHT;
		test_sprite[339] = WHT;
		test_sprite[340] = BLU;
		test_sprite[341] = BLU;
		test_sprite[342] = BLK;
		test_sprite[343] = BLK;
		test_sprite[344] = BLK;
		test_sprite[345] = BLK;
		test_sprite[346] = BLK;
		test_sprite[347] = BLK;
		test_sprite[348] = BLK;
		test_sprite[349] = BLK;
		test_sprite[350] = BLK;
		test_sprite[351] = BLK;
		test_sprite[352] = BLK;
		test_sprite[353] = BLK;
		test_sprite[354] = BLK;
		test_sprite[355] = BLK;
		test_sprite[356] = BLK;
		test_sprite[357] = BLK;
		test_sprite[358] = BLK;
		test_sprite[359] = BLK;
		test_sprite[360] = BLK;
		test_sprite[361] = RED;
		test_sprite[362] = RED;
		test_sprite[363] = RED;
		test_sprite[364] = WHT;
		test_sprite[365] = WHT;
		test_sprite[366] = BLU;
		test_sprite[367] = BLU;
		test_sprite[368] = RED;
		test_sprite[369] = RED;
		test_sprite[370] = WHT;
		test_sprite[371] = WHT;
		test_sprite[372] = BLU;
		test_sprite[373] = BLU;
		test_sprite[374] = RED;
		test_sprite[375] = BLK;
		test_sprite[376] = BLK;
		test_sprite[377] = BLK;
		test_sprite[378] = BLK;
		test_sprite[379] = BLK;
		test_sprite[380] = BLK;
		test_sprite[381] = BLK;
		test_sprite[382] = BLK;
		test_sprite[383] = BLK;
		test_sprite[384] = BLK;
		test_sprite[385] = BLK;
		test_sprite[386] = BLK;
		test_sprite[387] = BLK;
		test_sprite[388] = BLK;
		test_sprite[389] = BLK;
		test_sprite[390] = BLK;
		test_sprite[391] = BLK;
		test_sprite[392] = BLK;
		test_sprite[393] = RED;
		test_sprite[394] = RED;
		test_sprite[395] = RED;
		test_sprite[396] = RED;
		test_sprite[397] = WHT;
		test_sprite[398] = WHT;
		test_sprite[399] = RED;
		test_sprite[400] = RED;
		test_sprite[401] = RED;
		test_sprite[402] = RED;
		test_sprite[403] = WHT;
		test_sprite[404] = WHT;
		test_sprite[405] = RED;
		test_sprite[406] = RED;
		test_sprite[407] = BLK;
		test_sprite[408] = BLK;
		test_sprite[409] = BLK;
		test_sprite[410] = BLK;
		test_sprite[411] = BLK;
		test_sprite[412] = BLK;
		test_sprite[413] = BLK;
		test_sprite[414] = BLK;
		test_sprite[415] = BLK;
		test_sprite[416] = BLK;
		test_sprite[417] = BLK;
		test_sprite[418] = BLK;
		test_sprite[419] = BLK;
		test_sprite[420] = BLK;
		test_sprite[421] = BLK;
		test_sprite[422] = BLK;
		test_sprite[423] = BLK;
		test_sprite[424] = BLK;
		test_sprite[425] = RED;
		test_sprite[426] = RED;
		test_sprite[427] = RED;
		test_sprite[428] = RED;
		test_sprite[429] = RED;
		test_sprite[430] = RED;
		test_sprite[431] = RED;
		test_sprite[432] = RED;
		test_sprite[433] = RED;
		test_sprite[434] = RED;
		test_sprite[435] = RED;
		test_sprite[436] = RED;
		test_sprite[437] = RED;
		test_sprite[438] = RED;
		test_sprite[439] = BLK;
		test_sprite[440] = BLK;
		test_sprite[441] = BLK;
		test_sprite[442] = BLK;
		test_sprite[443] = BLK;
		test_sprite[444] = BLK;
		test_sprite[445] = BLK;
		test_sprite[446] = BLK;
		test_sprite[447] = BLK;
		test_sprite[448] = BLK;
		test_sprite[449] = BLK;
		test_sprite[450] = BLK;
		test_sprite[451] = BLK;
		test_sprite[452] = BLK;
		test_sprite[453] = BLK;
		test_sprite[454] = BLK;
		test_sprite[455] = BLK;
		test_sprite[456] = BLK;
		test_sprite[457] = RED;
		test_sprite[458] = RED;
		test_sprite[459] = RED;
		test_sprite[460] = RED;
		test_sprite[461] = RED;
		test_sprite[462] = RED;
		test_sprite[463] = RED;
		test_sprite[464] = RED;
		test_sprite[465] = RED;
		test_sprite[466] = RED;
		test_sprite[467] = RED;
		test_sprite[468] = RED;
		test_sprite[469] = RED;
		test_sprite[470] = RED;
		test_sprite[471] = BLK;
		test_sprite[472] = BLK;
		test_sprite[473] = BLK;
		test_sprite[474] = BLK;
		test_sprite[475] = BLK;
		test_sprite[476] = BLK;
		test_sprite[477] = BLK;
		test_sprite[478] = BLK;
		test_sprite[479] = BLK;
		test_sprite[480] = BLK;
		test_sprite[481] = BLK;
		test_sprite[482] = BLK;
		test_sprite[483] = BLK;
		test_sprite[484] = BLK;
		test_sprite[485] = BLK;
		test_sprite[486] = BLK;
		test_sprite[487] = BLK;
		test_sprite[488] = BLK;
		test_sprite[489] = RED;
		test_sprite[490] = RED;
		test_sprite[491] = RED;
		test_sprite[492] = RED;
		test_sprite[493] = RED;
		test_sprite[494] = RED;
		test_sprite[495] = RED;
		test_sprite[496] = RED;
		test_sprite[497] = RED;
		test_sprite[498] = RED;
		test_sprite[499] = RED;
		test_sprite[500] = RED;
		test_sprite[501] = RED;
		test_sprite[502] = RED;
		test_sprite[503] = BLK;
		test_sprite[504] = BLK;
		test_sprite[505] = BLK;
		test_sprite[506] = BLK;
		test_sprite[507] = BLK;
		test_sprite[508] = BLK;
		test_sprite[509] = BLK;
		test_sprite[510] = BLK;
		test_sprite[511] = BLK;
		test_sprite[512] = BLK;
		test_sprite[513] = BLK;
		test_sprite[514] = BLK;
		test_sprite[515] = BLK;
		test_sprite[516] = BLK;
		test_sprite[517] = BLK;
		test_sprite[518] = BLK;
		test_sprite[519] = BLK;
		test_sprite[520] = BLK;
		test_sprite[521] = RED;
		test_sprite[522] = RED;
		test_sprite[523] = RED;
		test_sprite[524] = RED;
		test_sprite[525] = RED;
		test_sprite[526] = RED;
		test_sprite[527] = RED;
		test_sprite[528] = RED;
		test_sprite[529] = RED;
		test_sprite[530] = RED;
		test_sprite[531] = RED;
		test_sprite[532] = RED;
		test_sprite[533] = RED;
		test_sprite[534] = RED;
		test_sprite[535] = BLK;
		test_sprite[536] = BLK;
		test_sprite[537] = BLK;
		test_sprite[538] = BLK;
		test_sprite[539] = BLK;
		test_sprite[540] = BLK;
		test_sprite[541] = BLK;
		test_sprite[542] = BLK;
		test_sprite[543] = BLK;
		test_sprite[544] = BLK;
		test_sprite[545] = BLK;
		test_sprite[546] = BLK;
		test_sprite[547] = BLK;
		test_sprite[548] = BLK;
		test_sprite[549] = BLK;
		test_sprite[550] = BLK;
		test_sprite[551] = BLK;
		test_sprite[552] = BLK;
		test_sprite[553] = RED;
		test_sprite[554] = RED;
		test_sprite[555] = BLK;
		test_sprite[556] = RED;
		test_sprite[557] = RED;
		test_sprite[558] = RED;
		test_sprite[559] = BLK;
		test_sprite[560] = BLK;
		test_sprite[561] = RED;
		test_sprite[562] = RED;
		test_sprite[563] = RED;
		test_sprite[564] = BLK;
		test_sprite[565] = RED;
		test_sprite[566] = RED;
		test_sprite[567] = BLK;
		test_sprite[568] = BLK;
		test_sprite[569] = BLK;
		test_sprite[570] = BLK;
		test_sprite[571] = BLK;
		test_sprite[572] = BLK;
		test_sprite[573] = BLK;
		test_sprite[574] = BLK;
		test_sprite[575] = BLK;
		test_sprite[576] = BLK;
		test_sprite[577] = BLK;
		test_sprite[578] = BLK;
		test_sprite[579] = BLK;
		test_sprite[580] = BLK;
		test_sprite[581] = BLK;
		test_sprite[582] = BLK;
		test_sprite[583] = BLK;
		test_sprite[584] = BLK;
		test_sprite[585] = RED;
		test_sprite[586] = BLK;
		test_sprite[587] = BLK;
		test_sprite[588] = BLK;
		test_sprite[589] = RED;
		test_sprite[590] = RED;
		test_sprite[591] = BLK;
		test_sprite[592] = BLK;
		test_sprite[593] = RED;
		test_sprite[594] = RED;
		test_sprite[595] = BLK;
		test_sprite[596] = BLK;
		test_sprite[597] = BLK;
		test_sprite[598] = RED;
		test_sprite[599] = BLK;
		test_sprite[600] = BLK;
		test_sprite[601] = BLK;
		test_sprite[602] = BLK;
		test_sprite[603] = BLK;
		test_sprite[604] = BLK;
		test_sprite[605] = BLK;
		test_sprite[606] = BLK;
		test_sprite[607] = BLK;
		test_sprite[608] = BLK;
		test_sprite[609] = BLK;
		test_sprite[610] = BLK;
		test_sprite[611] = BLK;
		test_sprite[612] = BLK;
		test_sprite[613] = BLK;
		test_sprite[614] = BLK;
		test_sprite[615] = BLK;
		test_sprite[616] = BLK;
		test_sprite[617] = BLK;
		test_sprite[618] = BLK;
		test_sprite[619] = BLK;
		test_sprite[620] = BLK;
		test_sprite[621] = BLK;
		test_sprite[622] = BLK;
		test_sprite[623] = BLK;
		test_sprite[624] = BLK;
		test_sprite[625] = BLK;
		test_sprite[626] = BLK;
		test_sprite[627] = BLK;
		test_sprite[628] = BLK;
		test_sprite[629] = BLK;
		test_sprite[630] = BLK;
		test_sprite[631] = BLK;
		test_sprite[632] = BLK;
		test_sprite[633] = BLK;
		test_sprite[634] = BLK;
		test_sprite[635] = BLK;
		test_sprite[636] = BLK;
		test_sprite[637] = BLK;
		test_sprite[638] = BLK;
		test_sprite[639] = BLK;
		test_sprite[640] = BLK;
		test_sprite[641] = BLK;
		test_sprite[642] = BLK;
		test_sprite[643] = BLK;
		test_sprite[644] = BLK;
		test_sprite[645] = BLK;
		test_sprite[646] = BLK;
		test_sprite[647] = BLK;
		test_sprite[648] = BLK;
		test_sprite[649] = BLK;
		test_sprite[650] = BLK;
		test_sprite[651] = BLK;
		test_sprite[652] = BLK;
		test_sprite[653] = BLK;
		test_sprite[654] = BLK;
		test_sprite[655] = BLK;
		test_sprite[656] = BLK;
		test_sprite[657] = BLK;
		test_sprite[658] = BLK;
		test_sprite[659] = BLK;
		test_sprite[660] = BLK;
		test_sprite[661] = BLK;
		test_sprite[662] = BLK;
		test_sprite[663] = BLK;
		test_sprite[664] = BLK;
		test_sprite[665] = BLK;
		test_sprite[666] = BLK;
		test_sprite[667] = BLK;
		test_sprite[668] = BLK;
		test_sprite[669] = BLK;
		test_sprite[670] = BLK;
		test_sprite[671] = BLK;
		test_sprite[672] = BLK;
		test_sprite[673] = BLK;
		test_sprite[674] = BLK;
		test_sprite[675] = BLK;
		test_sprite[676] = BLK;
		test_sprite[677] = BLK;
		test_sprite[678] = BLK;
		test_sprite[679] = BLK;
		test_sprite[680] = BLK;
		test_sprite[681] = BLK;
		test_sprite[682] = BLK;
		test_sprite[683] = BLK;
		test_sprite[684] = BLK;
		test_sprite[685] = BLK;
		test_sprite[686] = BLK;
		test_sprite[687] = BLK;
		test_sprite[688] = BLK;
		test_sprite[689] = BLK;
		test_sprite[690] = BLK;
		test_sprite[691] = BLK;
		test_sprite[692] = BLK;
		test_sprite[693] = BLK;
		test_sprite[694] = BLK;
		test_sprite[695] = BLK;
		test_sprite[696] = BLK;
		test_sprite[697] = BLK;
		test_sprite[698] = BLK;
		test_sprite[699] = BLK;
		test_sprite[700] = BLK;
		test_sprite[701] = BLK;
		test_sprite[702] = BLK;
		test_sprite[703] = BLK;
		test_sprite[704] = BLK;
		test_sprite[705] = BLK;
		test_sprite[706] = BLK;
		test_sprite[707] = BLK;
		test_sprite[708] = BLK;
		test_sprite[709] = BLK;
		test_sprite[710] = BLK;
		test_sprite[711] = BLK;
		test_sprite[712] = BLK;
		test_sprite[713] = BLK;
		test_sprite[714] = BLK;
		test_sprite[715] = BLK;
		test_sprite[716] = BLK;
		test_sprite[717] = BLK;
		test_sprite[718] = BLK;
		test_sprite[719] = BLK;
		test_sprite[720] = BLK;
		test_sprite[721] = BLK;
		test_sprite[722] = BLK;
		test_sprite[723] = BLK;
		test_sprite[724] = BLK;
		test_sprite[725] = BLK;
		test_sprite[726] = BLK;
		test_sprite[727] = BLK;
		test_sprite[728] = BLK;
		test_sprite[729] = BLK;
		test_sprite[730] = BLK;
		test_sprite[731] = BLK;
		test_sprite[732] = BLK;
		test_sprite[733] = BLK;
		test_sprite[734] = BLK;
		test_sprite[735] = BLK;
		test_sprite[736] = BLK;
		test_sprite[737] = BLK;
		test_sprite[738] = BLK;
		test_sprite[739] = BLK;
		test_sprite[740] = BLK;
		test_sprite[741] = BLK;
		test_sprite[742] = BLK;
		test_sprite[743] = BLK;
		test_sprite[744] = BLK;
		test_sprite[745] = BLK;
		test_sprite[746] = BLK;
		test_sprite[747] = BLK;
		test_sprite[748] = BLK;
		test_sprite[749] = BLK;
		test_sprite[750] = BLK;
		test_sprite[751] = BLK;
		test_sprite[752] = BLK;
		test_sprite[753] = BLK;
		test_sprite[754] = BLK;
		test_sprite[755] = BLK;
		test_sprite[756] = BLK;
		test_sprite[757] = BLK;
		test_sprite[758] = BLK;
		test_sprite[759] = BLK;
		test_sprite[760] = BLK;
		test_sprite[761] = BLK;
		test_sprite[762] = BLK;
		test_sprite[763] = BLK;
		test_sprite[764] = BLK;
		test_sprite[765] = BLK;
		test_sprite[766] = BLK;
		test_sprite[767] = BLK;
	end

endmodule
