`timescale 1ns / 1ns
module bin_to_bcd_tb;
	reg [6:0] number;
	wire [3:0] bcd0;
	wire [3:0] bcd1;
	bin_to_bcd dut(number, bcd0, bcd1);

	initial begin
		number=7'd0; #10;
		number=7'd1; #10;
		number=7'd2; #10;
		number=7'd3; #10;
		number=7'd4; #10;
		number=7'd5; #10;
		number=7'd6; #10;
		number=7'd7; #10;
		number=7'd8; #10;
		number=7'd9; #10;
		number=7'd10; #10;
		number=7'd11; #10;
		number=7'd12; #10;
		number=7'd13; #10;
		number=7'd14; #10;
		number=7'd15; #10;
		number=7'd16; #10;
		number=7'd17; #10;
		number=7'd18; #10;
		number=7'd19; #10;
		number=7'd20; #10;
		number=7'd21; #10;
		number=7'd22; #10;
		number=7'd23; #10;
		number=7'd24; #10;
		number=7'd25; #10;
		number=7'd26; #10;
		number=7'd27; #10;
		number=7'd28; #10;
		number=7'd29; #10;
		number=7'd30; #10;
		number=7'd31; #10;
		number=7'd32; #10;
		number=7'd33; #10;
		number=7'd34; #10;
		number=7'd35; #10;
		number=7'd36; #10;
		number=7'd37; #10;
		number=7'd38; #10;
		number=7'd39; #10;
		number=7'd40; #10;
		number=7'd41; #10;
		number=7'd42; #10;
		number=7'd43; #10;
		number=7'd44; #10;
		number=7'd45; #10;
		number=7'd46; #10;
		number=7'd47; #10;
		number=7'd48; #10;
		number=7'd49; #10;
		number=7'd50; #10;
		number=7'd51; #10;
		number=7'd52; #10;
		number=7'd53; #10;
		number=7'd54; #10;
		number=7'd55; #10;
		number=7'd56; #10;
		number=7'd57; #10;
		number=7'd58; #10;
		number=7'd59; #10;
		number=7'd60; #10;
		number=7'd61; #10;
		number=7'd62; #10;
		number=7'd63; #10;
		number=7'd64; #10;
		number=7'd65; #10;
		number=7'd66; #10;
		number=7'd67; #10;
		number=7'd68; #10;
		number=7'd69; #10;
		number=7'd70; #10;
		number=7'd71; #10;
		number=7'd72; #10;
		number=7'd73; #10;
		number=7'd74; #10;
		number=7'd75; #10;
		number=7'd76; #10;
		number=7'd77; #10;
		number=7'd78; #10;
		number=7'd79; #10;
		number=7'd80; #10;
		number=7'd81; #10;
		number=7'd82; #10;
		number=7'd83; #10;
		number=7'd84; #10;
		number=7'd85; #10;
		number=7'd86; #10;
		number=7'd87; #10;
		number=7'd88; #10;
		number=7'd89; #10;
		number=7'd90; #10;
		number=7'd91; #10;
		number=7'd92; #10;
		number=7'd93; #10;
		number=7'd94; #10;
		number=7'd95; #10;
		number=7'd96; #10;
		number=7'd97; #10;
		number=7'd98; #10;
		number=7'd99; #10;
	end

	initial begin
		$dumpfile("dump.vcd");
		$dumpvars();
	end
endmodule
