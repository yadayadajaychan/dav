module graphics(
	input vgaclk, // 25 MHz
	input rst, // active low

	input [3:0] grid [0:15],
	input [1:0] state,
	input [9:0] hc,
	input [9:0] vc,

	output reg [11:0] color // RGB
);

	reg bitmap [0:3071];
	reg [11:0] palette [0:23];

	reg [6:0] x;
	reg [6:0] y;
	assign x = hc/7;
	assign y = vc/7;

	reg [3:0] xi;
	reg [3:0] yi;
	assign xi = x % 16;
	assign yi = y % 16;

	reg [3:0] block;
	assign block = x/16 + y/4;

	always @(posedge vgaclk) begin
		if (x >= 64 || y >= 64 || block >= 16) begin
			color <= 12'd0;
		end else begin
			color <= palette[grid[block]*2 + bitmap[grid[block]*256 + xi + yi*16]];
		end
	end

	assign bitmap[0] = 1'b0;
	assign bitmap[1] = 1'b0;
	assign bitmap[2] = 1'b0;
	assign bitmap[3] = 1'b0;
	assign bitmap[4] = 1'b0;
	assign bitmap[5] = 1'b0;
	assign bitmap[6] = 1'b0;
	assign bitmap[7] = 1'b0;
	assign bitmap[8] = 1'b0;
	assign bitmap[9] = 1'b0;
	assign bitmap[10] = 1'b0;
	assign bitmap[11] = 1'b0;
	assign bitmap[12] = 1'b0;
	assign bitmap[13] = 1'b0;
	assign bitmap[14] = 1'b0;
	assign bitmap[15] = 1'b0;
	assign bitmap[16] = 1'b0;
	assign bitmap[17] = 1'b0;
	assign bitmap[18] = 1'b0;
	assign bitmap[19] = 1'b0;
	assign bitmap[20] = 1'b0;
	assign bitmap[21] = 1'b0;
	assign bitmap[22] = 1'b0;
	assign bitmap[23] = 1'b0;
	assign bitmap[24] = 1'b0;
	assign bitmap[25] = 1'b0;
	assign bitmap[26] = 1'b0;
	assign bitmap[27] = 1'b0;
	assign bitmap[28] = 1'b0;
	assign bitmap[29] = 1'b0;
	assign bitmap[30] = 1'b0;
	assign bitmap[31] = 1'b0;
	assign bitmap[32] = 1'b0;
	assign bitmap[33] = 1'b0;
	assign bitmap[34] = 1'b0;
	assign bitmap[35] = 1'b0;
	assign bitmap[36] = 1'b0;
	assign bitmap[37] = 1'b0;
	assign bitmap[38] = 1'b0;
	assign bitmap[39] = 1'b0;
	assign bitmap[40] = 1'b0;
	assign bitmap[41] = 1'b0;
	assign bitmap[42] = 1'b0;
	assign bitmap[43] = 1'b0;
	assign bitmap[44] = 1'b0;
	assign bitmap[45] = 1'b0;
	assign bitmap[46] = 1'b0;
	assign bitmap[47] = 1'b0;
	assign bitmap[48] = 1'b0;
	assign bitmap[49] = 1'b0;
	assign bitmap[50] = 1'b0;
	assign bitmap[51] = 1'b0;
	assign bitmap[52] = 1'b0;
	assign bitmap[53] = 1'b0;
	assign bitmap[54] = 1'b0;
	assign bitmap[55] = 1'b0;
	assign bitmap[56] = 1'b0;
	assign bitmap[57] = 1'b0;
	assign bitmap[58] = 1'b0;
	assign bitmap[59] = 1'b0;
	assign bitmap[60] = 1'b0;
	assign bitmap[61] = 1'b0;
	assign bitmap[62] = 1'b0;
	assign bitmap[63] = 1'b0;
	assign bitmap[64] = 1'b0;
	assign bitmap[65] = 1'b0;
	assign bitmap[66] = 1'b0;
	assign bitmap[67] = 1'b0;
	assign bitmap[68] = 1'b0;
	assign bitmap[69] = 1'b0;
	assign bitmap[70] = 1'b0;
	assign bitmap[71] = 1'b0;
	assign bitmap[72] = 1'b0;
	assign bitmap[73] = 1'b0;
	assign bitmap[74] = 1'b0;
	assign bitmap[75] = 1'b0;
	assign bitmap[76] = 1'b0;
	assign bitmap[77] = 1'b0;
	assign bitmap[78] = 1'b0;
	assign bitmap[79] = 1'b0;
	assign bitmap[80] = 1'b0;
	assign bitmap[81] = 1'b0;
	assign bitmap[82] = 1'b0;
	assign bitmap[83] = 1'b0;
	assign bitmap[84] = 1'b0;
	assign bitmap[85] = 1'b0;
	assign bitmap[86] = 1'b0;
	assign bitmap[87] = 1'b0;
	assign bitmap[88] = 1'b0;
	assign bitmap[89] = 1'b0;
	assign bitmap[90] = 1'b0;
	assign bitmap[91] = 1'b0;
	assign bitmap[92] = 1'b0;
	assign bitmap[93] = 1'b0;
	assign bitmap[94] = 1'b0;
	assign bitmap[95] = 1'b0;
	assign bitmap[96] = 1'b0;
	assign bitmap[97] = 1'b0;
	assign bitmap[98] = 1'b0;
	assign bitmap[99] = 1'b0;
	assign bitmap[100] = 1'b0;
	assign bitmap[101] = 1'b0;
	assign bitmap[102] = 1'b0;
	assign bitmap[103] = 1'b0;
	assign bitmap[104] = 1'b0;
	assign bitmap[105] = 1'b0;
	assign bitmap[106] = 1'b0;
	assign bitmap[107] = 1'b0;
	assign bitmap[108] = 1'b0;
	assign bitmap[109] = 1'b0;
	assign bitmap[110] = 1'b0;
	assign bitmap[111] = 1'b0;
	assign bitmap[112] = 1'b0;
	assign bitmap[113] = 1'b0;
	assign bitmap[114] = 1'b0;
	assign bitmap[115] = 1'b0;
	assign bitmap[116] = 1'b0;
	assign bitmap[117] = 1'b0;
	assign bitmap[118] = 1'b0;
	assign bitmap[119] = 1'b0;
	assign bitmap[120] = 1'b0;
	assign bitmap[121] = 1'b0;
	assign bitmap[122] = 1'b0;
	assign bitmap[123] = 1'b0;
	assign bitmap[124] = 1'b0;
	assign bitmap[125] = 1'b0;
	assign bitmap[126] = 1'b0;
	assign bitmap[127] = 1'b0;
	assign bitmap[128] = 1'b0;
	assign bitmap[129] = 1'b0;
	assign bitmap[130] = 1'b0;
	assign bitmap[131] = 1'b0;
	assign bitmap[132] = 1'b0;
	assign bitmap[133] = 1'b0;
	assign bitmap[134] = 1'b0;
	assign bitmap[135] = 1'b0;
	assign bitmap[136] = 1'b0;
	assign bitmap[137] = 1'b0;
	assign bitmap[138] = 1'b0;
	assign bitmap[139] = 1'b0;
	assign bitmap[140] = 1'b0;
	assign bitmap[141] = 1'b0;
	assign bitmap[142] = 1'b0;
	assign bitmap[143] = 1'b0;
	assign bitmap[144] = 1'b0;
	assign bitmap[145] = 1'b0;
	assign bitmap[146] = 1'b0;
	assign bitmap[147] = 1'b0;
	assign bitmap[148] = 1'b0;
	assign bitmap[149] = 1'b0;
	assign bitmap[150] = 1'b0;
	assign bitmap[151] = 1'b0;
	assign bitmap[152] = 1'b0;
	assign bitmap[153] = 1'b0;
	assign bitmap[154] = 1'b0;
	assign bitmap[155] = 1'b0;
	assign bitmap[156] = 1'b0;
	assign bitmap[157] = 1'b0;
	assign bitmap[158] = 1'b0;
	assign bitmap[159] = 1'b0;
	assign bitmap[160] = 1'b0;
	assign bitmap[161] = 1'b0;
	assign bitmap[162] = 1'b0;
	assign bitmap[163] = 1'b0;
	assign bitmap[164] = 1'b0;
	assign bitmap[165] = 1'b0;
	assign bitmap[166] = 1'b0;
	assign bitmap[167] = 1'b0;
	assign bitmap[168] = 1'b0;
	assign bitmap[169] = 1'b0;
	assign bitmap[170] = 1'b0;
	assign bitmap[171] = 1'b0;
	assign bitmap[172] = 1'b0;
	assign bitmap[173] = 1'b0;
	assign bitmap[174] = 1'b0;
	assign bitmap[175] = 1'b0;
	assign bitmap[176] = 1'b0;
	assign bitmap[177] = 1'b0;
	assign bitmap[178] = 1'b0;
	assign bitmap[179] = 1'b0;
	assign bitmap[180] = 1'b0;
	assign bitmap[181] = 1'b0;
	assign bitmap[182] = 1'b0;
	assign bitmap[183] = 1'b0;
	assign bitmap[184] = 1'b0;
	assign bitmap[185] = 1'b0;
	assign bitmap[186] = 1'b0;
	assign bitmap[187] = 1'b0;
	assign bitmap[188] = 1'b0;
	assign bitmap[189] = 1'b0;
	assign bitmap[190] = 1'b0;
	assign bitmap[191] = 1'b0;
	assign bitmap[192] = 1'b0;
	assign bitmap[193] = 1'b0;
	assign bitmap[194] = 1'b0;
	assign bitmap[195] = 1'b0;
	assign bitmap[196] = 1'b0;
	assign bitmap[197] = 1'b0;
	assign bitmap[198] = 1'b0;
	assign bitmap[199] = 1'b0;
	assign bitmap[200] = 1'b0;
	assign bitmap[201] = 1'b0;
	assign bitmap[202] = 1'b0;
	assign bitmap[203] = 1'b0;
	assign bitmap[204] = 1'b0;
	assign bitmap[205] = 1'b0;
	assign bitmap[206] = 1'b0;
	assign bitmap[207] = 1'b0;
	assign bitmap[208] = 1'b0;
	assign bitmap[209] = 1'b0;
	assign bitmap[210] = 1'b0;
	assign bitmap[211] = 1'b0;
	assign bitmap[212] = 1'b0;
	assign bitmap[213] = 1'b0;
	assign bitmap[214] = 1'b0;
	assign bitmap[215] = 1'b0;
	assign bitmap[216] = 1'b0;
	assign bitmap[217] = 1'b0;
	assign bitmap[218] = 1'b0;
	assign bitmap[219] = 1'b0;
	assign bitmap[220] = 1'b0;
	assign bitmap[221] = 1'b0;
	assign bitmap[222] = 1'b0;
	assign bitmap[223] = 1'b0;
	assign bitmap[224] = 1'b0;
	assign bitmap[225] = 1'b0;
	assign bitmap[226] = 1'b0;
	assign bitmap[227] = 1'b0;
	assign bitmap[228] = 1'b0;
	assign bitmap[229] = 1'b0;
	assign bitmap[230] = 1'b0;
	assign bitmap[231] = 1'b0;
	assign bitmap[232] = 1'b0;
	assign bitmap[233] = 1'b0;
	assign bitmap[234] = 1'b0;
	assign bitmap[235] = 1'b0;
	assign bitmap[236] = 1'b0;
	assign bitmap[237] = 1'b0;
	assign bitmap[238] = 1'b0;
	assign bitmap[239] = 1'b0;
	assign bitmap[240] = 1'b0;
	assign bitmap[241] = 1'b0;
	assign bitmap[242] = 1'b0;
	assign bitmap[243] = 1'b0;
	assign bitmap[244] = 1'b0;
	assign bitmap[245] = 1'b0;
	assign bitmap[246] = 1'b0;
	assign bitmap[247] = 1'b0;
	assign bitmap[248] = 1'b0;
	assign bitmap[249] = 1'b0;
	assign bitmap[250] = 1'b0;
	assign bitmap[251] = 1'b0;
	assign bitmap[252] = 1'b0;
	assign bitmap[253] = 1'b0;
	assign bitmap[254] = 1'b0;
	assign bitmap[255] = 1'b0;
	assign bitmap[256] = 1'b0;
	assign bitmap[257] = 1'b0;
	assign bitmap[258] = 1'b0;
	assign bitmap[259] = 1'b0;
	assign bitmap[260] = 1'b0;
	assign bitmap[261] = 1'b0;
	assign bitmap[262] = 1'b0;
	assign bitmap[263] = 1'b0;
	assign bitmap[264] = 1'b0;
	assign bitmap[265] = 1'b0;
	assign bitmap[266] = 1'b0;
	assign bitmap[267] = 1'b0;
	assign bitmap[268] = 1'b0;
	assign bitmap[269] = 1'b0;
	assign bitmap[270] = 1'b0;
	assign bitmap[271] = 1'b0;
	assign bitmap[272] = 1'b0;
	assign bitmap[273] = 1'b0;
	assign bitmap[274] = 1'b0;
	assign bitmap[275] = 1'b1;
	assign bitmap[276] = 1'b1;
	assign bitmap[277] = 1'b0;
	assign bitmap[278] = 1'b0;
	assign bitmap[279] = 1'b0;
	assign bitmap[280] = 1'b0;
	assign bitmap[281] = 1'b0;
	assign bitmap[282] = 1'b0;
	assign bitmap[283] = 1'b0;
	assign bitmap[284] = 1'b0;
	assign bitmap[285] = 1'b0;
	assign bitmap[286] = 1'b0;
	assign bitmap[287] = 1'b0;
	assign bitmap[288] = 1'b0;
	assign bitmap[289] = 1'b0;
	assign bitmap[290] = 1'b1;
	assign bitmap[291] = 1'b0;
	assign bitmap[292] = 1'b0;
	assign bitmap[293] = 1'b1;
	assign bitmap[294] = 1'b0;
	assign bitmap[295] = 1'b0;
	assign bitmap[296] = 1'b0;
	assign bitmap[297] = 1'b0;
	assign bitmap[298] = 1'b0;
	assign bitmap[299] = 1'b0;
	assign bitmap[300] = 1'b0;
	assign bitmap[301] = 1'b0;
	assign bitmap[302] = 1'b0;
	assign bitmap[303] = 1'b0;
	assign bitmap[304] = 1'b0;
	assign bitmap[305] = 1'b0;
	assign bitmap[306] = 1'b0;
	assign bitmap[307] = 1'b0;
	assign bitmap[308] = 1'b0;
	assign bitmap[309] = 1'b1;
	assign bitmap[310] = 1'b0;
	assign bitmap[311] = 1'b0;
	assign bitmap[312] = 1'b0;
	assign bitmap[313] = 1'b0;
	assign bitmap[314] = 1'b0;
	assign bitmap[315] = 1'b0;
	assign bitmap[316] = 1'b0;
	assign bitmap[317] = 1'b0;
	assign bitmap[318] = 1'b0;
	assign bitmap[319] = 1'b0;
	assign bitmap[320] = 1'b0;
	assign bitmap[321] = 1'b0;
	assign bitmap[322] = 1'b0;
	assign bitmap[323] = 1'b0;
	assign bitmap[324] = 1'b1;
	assign bitmap[325] = 1'b0;
	assign bitmap[326] = 1'b0;
	assign bitmap[327] = 1'b0;
	assign bitmap[328] = 1'b0;
	assign bitmap[329] = 1'b0;
	assign bitmap[330] = 1'b0;
	assign bitmap[331] = 1'b0;
	assign bitmap[332] = 1'b0;
	assign bitmap[333] = 1'b0;
	assign bitmap[334] = 1'b0;
	assign bitmap[335] = 1'b0;
	assign bitmap[336] = 1'b0;
	assign bitmap[337] = 1'b0;
	assign bitmap[338] = 1'b0;
	assign bitmap[339] = 1'b1;
	assign bitmap[340] = 1'b0;
	assign bitmap[341] = 1'b0;
	assign bitmap[342] = 1'b0;
	assign bitmap[343] = 1'b0;
	assign bitmap[344] = 1'b0;
	assign bitmap[345] = 1'b0;
	assign bitmap[346] = 1'b0;
	assign bitmap[347] = 1'b0;
	assign bitmap[348] = 1'b0;
	assign bitmap[349] = 1'b0;
	assign bitmap[350] = 1'b0;
	assign bitmap[351] = 1'b0;
	assign bitmap[352] = 1'b0;
	assign bitmap[353] = 1'b0;
	assign bitmap[354] = 1'b1;
	assign bitmap[355] = 1'b1;
	assign bitmap[356] = 1'b1;
	assign bitmap[357] = 1'b1;
	assign bitmap[358] = 1'b0;
	assign bitmap[359] = 1'b0;
	assign bitmap[360] = 1'b0;
	assign bitmap[361] = 1'b0;
	assign bitmap[362] = 1'b0;
	assign bitmap[363] = 1'b0;
	assign bitmap[364] = 1'b0;
	assign bitmap[365] = 1'b0;
	assign bitmap[366] = 1'b0;
	assign bitmap[367] = 1'b0;
	assign bitmap[368] = 1'b0;
	assign bitmap[369] = 1'b0;
	assign bitmap[370] = 1'b0;
	assign bitmap[371] = 1'b0;
	assign bitmap[372] = 1'b0;
	assign bitmap[373] = 1'b0;
	assign bitmap[374] = 1'b0;
	assign bitmap[375] = 1'b0;
	assign bitmap[376] = 1'b0;
	assign bitmap[377] = 1'b0;
	assign bitmap[378] = 1'b0;
	assign bitmap[379] = 1'b0;
	assign bitmap[380] = 1'b0;
	assign bitmap[381] = 1'b0;
	assign bitmap[382] = 1'b0;
	assign bitmap[383] = 1'b0;
	assign bitmap[384] = 1'b0;
	assign bitmap[385] = 1'b0;
	assign bitmap[386] = 1'b0;
	assign bitmap[387] = 1'b0;
	assign bitmap[388] = 1'b0;
	assign bitmap[389] = 1'b0;
	assign bitmap[390] = 1'b0;
	assign bitmap[391] = 1'b0;
	assign bitmap[392] = 1'b0;
	assign bitmap[393] = 1'b0;
	assign bitmap[394] = 1'b0;
	assign bitmap[395] = 1'b0;
	assign bitmap[396] = 1'b0;
	assign bitmap[397] = 1'b0;
	assign bitmap[398] = 1'b0;
	assign bitmap[399] = 1'b0;
	assign bitmap[400] = 1'b0;
	assign bitmap[401] = 1'b0;
	assign bitmap[402] = 1'b0;
	assign bitmap[403] = 1'b0;
	assign bitmap[404] = 1'b0;
	assign bitmap[405] = 1'b0;
	assign bitmap[406] = 1'b0;
	assign bitmap[407] = 1'b0;
	assign bitmap[408] = 1'b0;
	assign bitmap[409] = 1'b0;
	assign bitmap[410] = 1'b0;
	assign bitmap[411] = 1'b0;
	assign bitmap[412] = 1'b0;
	assign bitmap[413] = 1'b0;
	assign bitmap[414] = 1'b0;
	assign bitmap[415] = 1'b0;
	assign bitmap[416] = 1'b0;
	assign bitmap[417] = 1'b0;
	assign bitmap[418] = 1'b0;
	assign bitmap[419] = 1'b0;
	assign bitmap[420] = 1'b0;
	assign bitmap[421] = 1'b0;
	assign bitmap[422] = 1'b0;
	assign bitmap[423] = 1'b0;
	assign bitmap[424] = 1'b0;
	assign bitmap[425] = 1'b0;
	assign bitmap[426] = 1'b0;
	assign bitmap[427] = 1'b0;
	assign bitmap[428] = 1'b0;
	assign bitmap[429] = 1'b0;
	assign bitmap[430] = 1'b0;
	assign bitmap[431] = 1'b0;
	assign bitmap[432] = 1'b0;
	assign bitmap[433] = 1'b0;
	assign bitmap[434] = 1'b0;
	assign bitmap[435] = 1'b0;
	assign bitmap[436] = 1'b0;
	assign bitmap[437] = 1'b0;
	assign bitmap[438] = 1'b0;
	assign bitmap[439] = 1'b0;
	assign bitmap[440] = 1'b0;
	assign bitmap[441] = 1'b0;
	assign bitmap[442] = 1'b0;
	assign bitmap[443] = 1'b0;
	assign bitmap[444] = 1'b0;
	assign bitmap[445] = 1'b0;
	assign bitmap[446] = 1'b0;
	assign bitmap[447] = 1'b0;
	assign bitmap[448] = 1'b0;
	assign bitmap[449] = 1'b0;
	assign bitmap[450] = 1'b0;
	assign bitmap[451] = 1'b0;
	assign bitmap[452] = 1'b0;
	assign bitmap[453] = 1'b0;
	assign bitmap[454] = 1'b0;
	assign bitmap[455] = 1'b0;
	assign bitmap[456] = 1'b0;
	assign bitmap[457] = 1'b0;
	assign bitmap[458] = 1'b0;
	assign bitmap[459] = 1'b0;
	assign bitmap[460] = 1'b0;
	assign bitmap[461] = 1'b0;
	assign bitmap[462] = 1'b0;
	assign bitmap[463] = 1'b0;
	assign bitmap[464] = 1'b0;
	assign bitmap[465] = 1'b0;
	assign bitmap[466] = 1'b0;
	assign bitmap[467] = 1'b0;
	assign bitmap[468] = 1'b0;
	assign bitmap[469] = 1'b0;
	assign bitmap[470] = 1'b0;
	assign bitmap[471] = 1'b0;
	assign bitmap[472] = 1'b0;
	assign bitmap[473] = 1'b0;
	assign bitmap[474] = 1'b0;
	assign bitmap[475] = 1'b0;
	assign bitmap[476] = 1'b0;
	assign bitmap[477] = 1'b0;
	assign bitmap[478] = 1'b0;
	assign bitmap[479] = 1'b0;
	assign bitmap[480] = 1'b0;
	assign bitmap[481] = 1'b0;
	assign bitmap[482] = 1'b0;
	assign bitmap[483] = 1'b0;
	assign bitmap[484] = 1'b0;
	assign bitmap[485] = 1'b0;
	assign bitmap[486] = 1'b0;
	assign bitmap[487] = 1'b0;
	assign bitmap[488] = 1'b0;
	assign bitmap[489] = 1'b0;
	assign bitmap[490] = 1'b0;
	assign bitmap[491] = 1'b0;
	assign bitmap[492] = 1'b0;
	assign bitmap[493] = 1'b0;
	assign bitmap[494] = 1'b0;
	assign bitmap[495] = 1'b0;
	assign bitmap[496] = 1'b0;
	assign bitmap[497] = 1'b0;
	assign bitmap[498] = 1'b0;
	assign bitmap[499] = 1'b0;
	assign bitmap[500] = 1'b0;
	assign bitmap[501] = 1'b0;
	assign bitmap[502] = 1'b0;
	assign bitmap[503] = 1'b0;
	assign bitmap[504] = 1'b0;
	assign bitmap[505] = 1'b0;
	assign bitmap[506] = 1'b0;
	assign bitmap[507] = 1'b0;
	assign bitmap[508] = 1'b0;
	assign bitmap[509] = 1'b0;
	assign bitmap[510] = 1'b0;
	assign bitmap[511] = 1'b0;
	assign bitmap[512] = 1'b0;
	assign bitmap[513] = 1'b0;
	assign bitmap[514] = 1'b0;
	assign bitmap[515] = 1'b0;
	assign bitmap[516] = 1'b0;
	assign bitmap[517] = 1'b0;
	assign bitmap[518] = 1'b0;
	assign bitmap[519] = 1'b0;
	assign bitmap[520] = 1'b0;
	assign bitmap[521] = 1'b0;
	assign bitmap[522] = 1'b0;
	assign bitmap[523] = 1'b0;
	assign bitmap[524] = 1'b0;
	assign bitmap[525] = 1'b0;
	assign bitmap[526] = 1'b0;
	assign bitmap[527] = 1'b0;
	assign bitmap[528] = 1'b0;
	assign bitmap[529] = 1'b0;
	assign bitmap[530] = 1'b0;
	assign bitmap[531] = 1'b0;
	assign bitmap[532] = 1'b1;
	assign bitmap[533] = 1'b1;
	assign bitmap[534] = 1'b0;
	assign bitmap[535] = 1'b0;
	assign bitmap[536] = 1'b0;
	assign bitmap[537] = 1'b0;
	assign bitmap[538] = 1'b0;
	assign bitmap[539] = 1'b0;
	assign bitmap[540] = 1'b0;
	assign bitmap[541] = 1'b0;
	assign bitmap[542] = 1'b0;
	assign bitmap[543] = 1'b0;
	assign bitmap[544] = 1'b0;
	assign bitmap[545] = 1'b0;
	assign bitmap[546] = 1'b0;
	assign bitmap[547] = 1'b1;
	assign bitmap[548] = 1'b0;
	assign bitmap[549] = 1'b1;
	assign bitmap[550] = 1'b0;
	assign bitmap[551] = 1'b0;
	assign bitmap[552] = 1'b0;
	assign bitmap[553] = 1'b0;
	assign bitmap[554] = 1'b0;
	assign bitmap[555] = 1'b0;
	assign bitmap[556] = 1'b0;
	assign bitmap[557] = 1'b0;
	assign bitmap[558] = 1'b0;
	assign bitmap[559] = 1'b0;
	assign bitmap[560] = 1'b0;
	assign bitmap[561] = 1'b0;
	assign bitmap[562] = 1'b1;
	assign bitmap[563] = 1'b0;
	assign bitmap[564] = 1'b0;
	assign bitmap[565] = 1'b1;
	assign bitmap[566] = 1'b0;
	assign bitmap[567] = 1'b0;
	assign bitmap[568] = 1'b0;
	assign bitmap[569] = 1'b0;
	assign bitmap[570] = 1'b0;
	assign bitmap[571] = 1'b0;
	assign bitmap[572] = 1'b0;
	assign bitmap[573] = 1'b0;
	assign bitmap[574] = 1'b0;
	assign bitmap[575] = 1'b0;
	assign bitmap[576] = 1'b0;
	assign bitmap[577] = 1'b0;
	assign bitmap[578] = 1'b1;
	assign bitmap[579] = 1'b1;
	assign bitmap[580] = 1'b1;
	assign bitmap[581] = 1'b1;
	assign bitmap[582] = 1'b1;
	assign bitmap[583] = 1'b0;
	assign bitmap[584] = 1'b0;
	assign bitmap[585] = 1'b0;
	assign bitmap[586] = 1'b0;
	assign bitmap[587] = 1'b0;
	assign bitmap[588] = 1'b0;
	assign bitmap[589] = 1'b0;
	assign bitmap[590] = 1'b0;
	assign bitmap[591] = 1'b0;
	assign bitmap[592] = 1'b0;
	assign bitmap[593] = 1'b0;
	assign bitmap[594] = 1'b0;
	assign bitmap[595] = 1'b0;
	assign bitmap[596] = 1'b0;
	assign bitmap[597] = 1'b1;
	assign bitmap[598] = 1'b0;
	assign bitmap[599] = 1'b0;
	assign bitmap[600] = 1'b0;
	assign bitmap[601] = 1'b0;
	assign bitmap[602] = 1'b0;
	assign bitmap[603] = 1'b0;
	assign bitmap[604] = 1'b0;
	assign bitmap[605] = 1'b0;
	assign bitmap[606] = 1'b0;
	assign bitmap[607] = 1'b0;
	assign bitmap[608] = 1'b0;
	assign bitmap[609] = 1'b0;
	assign bitmap[610] = 1'b0;
	assign bitmap[611] = 1'b0;
	assign bitmap[612] = 1'b0;
	assign bitmap[613] = 1'b1;
	assign bitmap[614] = 1'b0;
	assign bitmap[615] = 1'b0;
	assign bitmap[616] = 1'b0;
	assign bitmap[617] = 1'b0;
	assign bitmap[618] = 1'b0;
	assign bitmap[619] = 1'b0;
	assign bitmap[620] = 1'b0;
	assign bitmap[621] = 1'b0;
	assign bitmap[622] = 1'b0;
	assign bitmap[623] = 1'b0;
	assign bitmap[624] = 1'b0;
	assign bitmap[625] = 1'b0;
	assign bitmap[626] = 1'b0;
	assign bitmap[627] = 1'b0;
	assign bitmap[628] = 1'b0;
	assign bitmap[629] = 1'b0;
	assign bitmap[630] = 1'b0;
	assign bitmap[631] = 1'b0;
	assign bitmap[632] = 1'b0;
	assign bitmap[633] = 1'b0;
	assign bitmap[634] = 1'b0;
	assign bitmap[635] = 1'b0;
	assign bitmap[636] = 1'b0;
	assign bitmap[637] = 1'b0;
	assign bitmap[638] = 1'b0;
	assign bitmap[639] = 1'b0;
	assign bitmap[640] = 1'b0;
	assign bitmap[641] = 1'b0;
	assign bitmap[642] = 1'b0;
	assign bitmap[643] = 1'b0;
	assign bitmap[644] = 1'b0;
	assign bitmap[645] = 1'b0;
	assign bitmap[646] = 1'b0;
	assign bitmap[647] = 1'b0;
	assign bitmap[648] = 1'b0;
	assign bitmap[649] = 1'b0;
	assign bitmap[650] = 1'b0;
	assign bitmap[651] = 1'b0;
	assign bitmap[652] = 1'b0;
	assign bitmap[653] = 1'b0;
	assign bitmap[654] = 1'b0;
	assign bitmap[655] = 1'b0;
	assign bitmap[656] = 1'b0;
	assign bitmap[657] = 1'b0;
	assign bitmap[658] = 1'b0;
	assign bitmap[659] = 1'b0;
	assign bitmap[660] = 1'b0;
	assign bitmap[661] = 1'b0;
	assign bitmap[662] = 1'b0;
	assign bitmap[663] = 1'b0;
	assign bitmap[664] = 1'b0;
	assign bitmap[665] = 1'b0;
	assign bitmap[666] = 1'b0;
	assign bitmap[667] = 1'b0;
	assign bitmap[668] = 1'b0;
	assign bitmap[669] = 1'b0;
	assign bitmap[670] = 1'b0;
	assign bitmap[671] = 1'b0;
	assign bitmap[672] = 1'b0;
	assign bitmap[673] = 1'b0;
	assign bitmap[674] = 1'b0;
	assign bitmap[675] = 1'b0;
	assign bitmap[676] = 1'b0;
	assign bitmap[677] = 1'b0;
	assign bitmap[678] = 1'b0;
	assign bitmap[679] = 1'b0;
	assign bitmap[680] = 1'b0;
	assign bitmap[681] = 1'b0;
	assign bitmap[682] = 1'b0;
	assign bitmap[683] = 1'b0;
	assign bitmap[684] = 1'b0;
	assign bitmap[685] = 1'b0;
	assign bitmap[686] = 1'b0;
	assign bitmap[687] = 1'b0;
	assign bitmap[688] = 1'b0;
	assign bitmap[689] = 1'b0;
	assign bitmap[690] = 1'b0;
	assign bitmap[691] = 1'b0;
	assign bitmap[692] = 1'b0;
	assign bitmap[693] = 1'b0;
	assign bitmap[694] = 1'b0;
	assign bitmap[695] = 1'b0;
	assign bitmap[696] = 1'b0;
	assign bitmap[697] = 1'b0;
	assign bitmap[698] = 1'b0;
	assign bitmap[699] = 1'b0;
	assign bitmap[700] = 1'b0;
	assign bitmap[701] = 1'b0;
	assign bitmap[702] = 1'b0;
	assign bitmap[703] = 1'b0;
	assign bitmap[704] = 1'b0;
	assign bitmap[705] = 1'b0;
	assign bitmap[706] = 1'b0;
	assign bitmap[707] = 1'b0;
	assign bitmap[708] = 1'b0;
	assign bitmap[709] = 1'b0;
	assign bitmap[710] = 1'b0;
	assign bitmap[711] = 1'b0;
	assign bitmap[712] = 1'b0;
	assign bitmap[713] = 1'b0;
	assign bitmap[714] = 1'b0;
	assign bitmap[715] = 1'b0;
	assign bitmap[716] = 1'b0;
	assign bitmap[717] = 1'b0;
	assign bitmap[718] = 1'b0;
	assign bitmap[719] = 1'b0;
	assign bitmap[720] = 1'b0;
	assign bitmap[721] = 1'b0;
	assign bitmap[722] = 1'b0;
	assign bitmap[723] = 1'b0;
	assign bitmap[724] = 1'b0;
	assign bitmap[725] = 1'b0;
	assign bitmap[726] = 1'b0;
	assign bitmap[727] = 1'b0;
	assign bitmap[728] = 1'b0;
	assign bitmap[729] = 1'b0;
	assign bitmap[730] = 1'b0;
	assign bitmap[731] = 1'b0;
	assign bitmap[732] = 1'b0;
	assign bitmap[733] = 1'b0;
	assign bitmap[734] = 1'b0;
	assign bitmap[735] = 1'b0;
	assign bitmap[736] = 1'b0;
	assign bitmap[737] = 1'b0;
	assign bitmap[738] = 1'b0;
	assign bitmap[739] = 1'b0;
	assign bitmap[740] = 1'b0;
	assign bitmap[741] = 1'b0;
	assign bitmap[742] = 1'b0;
	assign bitmap[743] = 1'b0;
	assign bitmap[744] = 1'b0;
	assign bitmap[745] = 1'b0;
	assign bitmap[746] = 1'b0;
	assign bitmap[747] = 1'b0;
	assign bitmap[748] = 1'b0;
	assign bitmap[749] = 1'b0;
	assign bitmap[750] = 1'b0;
	assign bitmap[751] = 1'b0;
	assign bitmap[752] = 1'b0;
	assign bitmap[753] = 1'b0;
	assign bitmap[754] = 1'b0;
	assign bitmap[755] = 1'b0;
	assign bitmap[756] = 1'b0;
	assign bitmap[757] = 1'b0;
	assign bitmap[758] = 1'b0;
	assign bitmap[759] = 1'b0;
	assign bitmap[760] = 1'b0;
	assign bitmap[761] = 1'b0;
	assign bitmap[762] = 1'b0;
	assign bitmap[763] = 1'b0;
	assign bitmap[764] = 1'b0;
	assign bitmap[765] = 1'b0;
	assign bitmap[766] = 1'b0;
	assign bitmap[767] = 1'b0;
	assign bitmap[768] = 1'b0;
	assign bitmap[769] = 1'b0;
	assign bitmap[770] = 1'b0;
	assign bitmap[771] = 1'b0;
	assign bitmap[772] = 1'b0;
	assign bitmap[773] = 1'b0;
	assign bitmap[774] = 1'b0;
	assign bitmap[775] = 1'b0;
	assign bitmap[776] = 1'b0;
	assign bitmap[777] = 1'b0;
	assign bitmap[778] = 1'b0;
	assign bitmap[779] = 1'b0;
	assign bitmap[780] = 1'b0;
	assign bitmap[781] = 1'b0;
	assign bitmap[782] = 1'b0;
	assign bitmap[783] = 1'b0;
	assign bitmap[784] = 1'b0;
	assign bitmap[785] = 1'b0;
	assign bitmap[786] = 1'b1;
	assign bitmap[787] = 1'b1;
	assign bitmap[788] = 1'b1;
	assign bitmap[789] = 1'b1;
	assign bitmap[790] = 1'b0;
	assign bitmap[791] = 1'b0;
	assign bitmap[792] = 1'b0;
	assign bitmap[793] = 1'b0;
	assign bitmap[794] = 1'b0;
	assign bitmap[795] = 1'b0;
	assign bitmap[796] = 1'b0;
	assign bitmap[797] = 1'b0;
	assign bitmap[798] = 1'b0;
	assign bitmap[799] = 1'b0;
	assign bitmap[800] = 1'b0;
	assign bitmap[801] = 1'b0;
	assign bitmap[802] = 1'b1;
	assign bitmap[803] = 1'b0;
	assign bitmap[804] = 1'b0;
	assign bitmap[805] = 1'b1;
	assign bitmap[806] = 1'b0;
	assign bitmap[807] = 1'b0;
	assign bitmap[808] = 1'b0;
	assign bitmap[809] = 1'b0;
	assign bitmap[810] = 1'b0;
	assign bitmap[811] = 1'b0;
	assign bitmap[812] = 1'b0;
	assign bitmap[813] = 1'b0;
	assign bitmap[814] = 1'b0;
	assign bitmap[815] = 1'b0;
	assign bitmap[816] = 1'b0;
	assign bitmap[817] = 1'b0;
	assign bitmap[818] = 1'b1;
	assign bitmap[819] = 1'b0;
	assign bitmap[820] = 1'b0;
	assign bitmap[821] = 1'b1;
	assign bitmap[822] = 1'b0;
	assign bitmap[823] = 1'b0;
	assign bitmap[824] = 1'b0;
	assign bitmap[825] = 1'b0;
	assign bitmap[826] = 1'b0;
	assign bitmap[827] = 1'b0;
	assign bitmap[828] = 1'b0;
	assign bitmap[829] = 1'b0;
	assign bitmap[830] = 1'b0;
	assign bitmap[831] = 1'b0;
	assign bitmap[832] = 1'b0;
	assign bitmap[833] = 1'b0;
	assign bitmap[834] = 1'b1;
	assign bitmap[835] = 1'b1;
	assign bitmap[836] = 1'b1;
	assign bitmap[837] = 1'b1;
	assign bitmap[838] = 1'b0;
	assign bitmap[839] = 1'b0;
	assign bitmap[840] = 1'b0;
	assign bitmap[841] = 1'b0;
	assign bitmap[842] = 1'b0;
	assign bitmap[843] = 1'b0;
	assign bitmap[844] = 1'b0;
	assign bitmap[845] = 1'b0;
	assign bitmap[846] = 1'b0;
	assign bitmap[847] = 1'b0;
	assign bitmap[848] = 1'b0;
	assign bitmap[849] = 1'b0;
	assign bitmap[850] = 1'b1;
	assign bitmap[851] = 1'b0;
	assign bitmap[852] = 1'b0;
	assign bitmap[853] = 1'b1;
	assign bitmap[854] = 1'b0;
	assign bitmap[855] = 1'b0;
	assign bitmap[856] = 1'b0;
	assign bitmap[857] = 1'b0;
	assign bitmap[858] = 1'b0;
	assign bitmap[859] = 1'b0;
	assign bitmap[860] = 1'b0;
	assign bitmap[861] = 1'b0;
	assign bitmap[862] = 1'b0;
	assign bitmap[863] = 1'b0;
	assign bitmap[864] = 1'b0;
	assign bitmap[865] = 1'b0;
	assign bitmap[866] = 1'b1;
	assign bitmap[867] = 1'b1;
	assign bitmap[868] = 1'b1;
	assign bitmap[869] = 1'b1;
	assign bitmap[870] = 1'b0;
	assign bitmap[871] = 1'b0;
	assign bitmap[872] = 1'b0;
	assign bitmap[873] = 1'b0;
	assign bitmap[874] = 1'b0;
	assign bitmap[875] = 1'b0;
	assign bitmap[876] = 1'b0;
	assign bitmap[877] = 1'b0;
	assign bitmap[878] = 1'b0;
	assign bitmap[879] = 1'b0;
	assign bitmap[880] = 1'b0;
	assign bitmap[881] = 1'b0;
	assign bitmap[882] = 1'b0;
	assign bitmap[883] = 1'b0;
	assign bitmap[884] = 1'b0;
	assign bitmap[885] = 1'b0;
	assign bitmap[886] = 1'b0;
	assign bitmap[887] = 1'b0;
	assign bitmap[888] = 1'b0;
	assign bitmap[889] = 1'b0;
	assign bitmap[890] = 1'b0;
	assign bitmap[891] = 1'b0;
	assign bitmap[892] = 1'b0;
	assign bitmap[893] = 1'b0;
	assign bitmap[894] = 1'b0;
	assign bitmap[895] = 1'b0;
	assign bitmap[896] = 1'b0;
	assign bitmap[897] = 1'b0;
	assign bitmap[898] = 1'b0;
	assign bitmap[899] = 1'b0;
	assign bitmap[900] = 1'b0;
	assign bitmap[901] = 1'b0;
	assign bitmap[902] = 1'b0;
	assign bitmap[903] = 1'b0;
	assign bitmap[904] = 1'b0;
	assign bitmap[905] = 1'b0;
	assign bitmap[906] = 1'b0;
	assign bitmap[907] = 1'b0;
	assign bitmap[908] = 1'b0;
	assign bitmap[909] = 1'b0;
	assign bitmap[910] = 1'b0;
	assign bitmap[911] = 1'b0;
	assign bitmap[912] = 1'b0;
	assign bitmap[913] = 1'b0;
	assign bitmap[914] = 1'b0;
	assign bitmap[915] = 1'b0;
	assign bitmap[916] = 1'b0;
	assign bitmap[917] = 1'b0;
	assign bitmap[918] = 1'b0;
	assign bitmap[919] = 1'b0;
	assign bitmap[920] = 1'b0;
	assign bitmap[921] = 1'b0;
	assign bitmap[922] = 1'b0;
	assign bitmap[923] = 1'b0;
	assign bitmap[924] = 1'b0;
	assign bitmap[925] = 1'b0;
	assign bitmap[926] = 1'b0;
	assign bitmap[927] = 1'b0;
	assign bitmap[928] = 1'b0;
	assign bitmap[929] = 1'b0;
	assign bitmap[930] = 1'b0;
	assign bitmap[931] = 1'b0;
	assign bitmap[932] = 1'b0;
	assign bitmap[933] = 1'b0;
	assign bitmap[934] = 1'b0;
	assign bitmap[935] = 1'b0;
	assign bitmap[936] = 1'b0;
	assign bitmap[937] = 1'b0;
	assign bitmap[938] = 1'b0;
	assign bitmap[939] = 1'b0;
	assign bitmap[940] = 1'b0;
	assign bitmap[941] = 1'b0;
	assign bitmap[942] = 1'b0;
	assign bitmap[943] = 1'b0;
	assign bitmap[944] = 1'b0;
	assign bitmap[945] = 1'b0;
	assign bitmap[946] = 1'b0;
	assign bitmap[947] = 1'b0;
	assign bitmap[948] = 1'b0;
	assign bitmap[949] = 1'b0;
	assign bitmap[950] = 1'b0;
	assign bitmap[951] = 1'b0;
	assign bitmap[952] = 1'b0;
	assign bitmap[953] = 1'b0;
	assign bitmap[954] = 1'b0;
	assign bitmap[955] = 1'b0;
	assign bitmap[956] = 1'b0;
	assign bitmap[957] = 1'b0;
	assign bitmap[958] = 1'b0;
	assign bitmap[959] = 1'b0;
	assign bitmap[960] = 1'b0;
	assign bitmap[961] = 1'b0;
	assign bitmap[962] = 1'b0;
	assign bitmap[963] = 1'b0;
	assign bitmap[964] = 1'b0;
	assign bitmap[965] = 1'b0;
	assign bitmap[966] = 1'b0;
	assign bitmap[967] = 1'b0;
	assign bitmap[968] = 1'b0;
	assign bitmap[969] = 1'b0;
	assign bitmap[970] = 1'b0;
	assign bitmap[971] = 1'b0;
	assign bitmap[972] = 1'b0;
	assign bitmap[973] = 1'b0;
	assign bitmap[974] = 1'b0;
	assign bitmap[975] = 1'b0;
	assign bitmap[976] = 1'b0;
	assign bitmap[977] = 1'b0;
	assign bitmap[978] = 1'b0;
	assign bitmap[979] = 1'b0;
	assign bitmap[980] = 1'b0;
	assign bitmap[981] = 1'b0;
	assign bitmap[982] = 1'b0;
	assign bitmap[983] = 1'b0;
	assign bitmap[984] = 1'b0;
	assign bitmap[985] = 1'b0;
	assign bitmap[986] = 1'b0;
	assign bitmap[987] = 1'b0;
	assign bitmap[988] = 1'b0;
	assign bitmap[989] = 1'b0;
	assign bitmap[990] = 1'b0;
	assign bitmap[991] = 1'b0;
	assign bitmap[992] = 1'b0;
	assign bitmap[993] = 1'b0;
	assign bitmap[994] = 1'b0;
	assign bitmap[995] = 1'b0;
	assign bitmap[996] = 1'b0;
	assign bitmap[997] = 1'b0;
	assign bitmap[998] = 1'b0;
	assign bitmap[999] = 1'b0;
	assign bitmap[1000] = 1'b0;
	assign bitmap[1001] = 1'b0;
	assign bitmap[1002] = 1'b0;
	assign bitmap[1003] = 1'b0;
	assign bitmap[1004] = 1'b0;
	assign bitmap[1005] = 1'b0;
	assign bitmap[1006] = 1'b0;
	assign bitmap[1007] = 1'b0;
	assign bitmap[1008] = 1'b0;
	assign bitmap[1009] = 1'b0;
	assign bitmap[1010] = 1'b0;
	assign bitmap[1011] = 1'b0;
	assign bitmap[1012] = 1'b0;
	assign bitmap[1013] = 1'b0;
	assign bitmap[1014] = 1'b0;
	assign bitmap[1015] = 1'b0;
	assign bitmap[1016] = 1'b0;
	assign bitmap[1017] = 1'b0;
	assign bitmap[1018] = 1'b0;
	assign bitmap[1019] = 1'b0;
	assign bitmap[1020] = 1'b0;
	assign bitmap[1021] = 1'b0;
	assign bitmap[1022] = 1'b0;
	assign bitmap[1023] = 1'b0;
	assign bitmap[1024] = 1'b0;
	assign bitmap[1025] = 1'b0;
	assign bitmap[1026] = 1'b0;
	assign bitmap[1027] = 1'b0;
	assign bitmap[1028] = 1'b0;
	assign bitmap[1029] = 1'b0;
	assign bitmap[1030] = 1'b0;
	assign bitmap[1031] = 1'b0;
	assign bitmap[1032] = 1'b0;
	assign bitmap[1033] = 1'b0;
	assign bitmap[1034] = 1'b0;
	assign bitmap[1035] = 1'b0;
	assign bitmap[1036] = 1'b0;
	assign bitmap[1037] = 1'b0;
	assign bitmap[1038] = 1'b0;
	assign bitmap[1039] = 1'b0;
	assign bitmap[1040] = 1'b0;
	assign bitmap[1041] = 1'b0;
	assign bitmap[1042] = 1'b0;
	assign bitmap[1043] = 1'b0;
	assign bitmap[1044] = 1'b1;
	assign bitmap[1045] = 1'b0;
	assign bitmap[1046] = 1'b0;
	assign bitmap[1047] = 1'b0;
	assign bitmap[1048] = 1'b0;
	assign bitmap[1049] = 1'b0;
	assign bitmap[1050] = 1'b1;
	assign bitmap[1051] = 1'b1;
	assign bitmap[1052] = 1'b1;
	assign bitmap[1053] = 1'b1;
	assign bitmap[1054] = 1'b0;
	assign bitmap[1055] = 1'b0;
	assign bitmap[1056] = 1'b0;
	assign bitmap[1057] = 1'b0;
	assign bitmap[1058] = 1'b0;
	assign bitmap[1059] = 1'b1;
	assign bitmap[1060] = 1'b1;
	assign bitmap[1061] = 1'b0;
	assign bitmap[1062] = 1'b0;
	assign bitmap[1063] = 1'b0;
	assign bitmap[1064] = 1'b0;
	assign bitmap[1065] = 1'b0;
	assign bitmap[1066] = 1'b1;
	assign bitmap[1067] = 1'b0;
	assign bitmap[1068] = 1'b0;
	assign bitmap[1069] = 1'b0;
	assign bitmap[1070] = 1'b0;
	assign bitmap[1071] = 1'b0;
	assign bitmap[1072] = 1'b0;
	assign bitmap[1073] = 1'b0;
	assign bitmap[1074] = 1'b1;
	assign bitmap[1075] = 1'b0;
	assign bitmap[1076] = 1'b1;
	assign bitmap[1077] = 1'b0;
	assign bitmap[1078] = 1'b0;
	assign bitmap[1079] = 1'b0;
	assign bitmap[1080] = 1'b0;
	assign bitmap[1081] = 1'b0;
	assign bitmap[1082] = 1'b1;
	assign bitmap[1083] = 1'b0;
	assign bitmap[1084] = 1'b0;
	assign bitmap[1085] = 1'b0;
	assign bitmap[1086] = 1'b0;
	assign bitmap[1087] = 1'b0;
	assign bitmap[1088] = 1'b0;
	assign bitmap[1089] = 1'b0;
	assign bitmap[1090] = 1'b0;
	assign bitmap[1091] = 1'b0;
	assign bitmap[1092] = 1'b1;
	assign bitmap[1093] = 1'b0;
	assign bitmap[1094] = 1'b0;
	assign bitmap[1095] = 1'b0;
	assign bitmap[1096] = 1'b0;
	assign bitmap[1097] = 1'b0;
	assign bitmap[1098] = 1'b1;
	assign bitmap[1099] = 1'b1;
	assign bitmap[1100] = 1'b1;
	assign bitmap[1101] = 1'b1;
	assign bitmap[1102] = 1'b0;
	assign bitmap[1103] = 1'b0;
	assign bitmap[1104] = 1'b0;
	assign bitmap[1105] = 1'b0;
	assign bitmap[1106] = 1'b0;
	assign bitmap[1107] = 1'b0;
	assign bitmap[1108] = 1'b1;
	assign bitmap[1109] = 1'b0;
	assign bitmap[1110] = 1'b0;
	assign bitmap[1111] = 1'b0;
	assign bitmap[1112] = 1'b0;
	assign bitmap[1113] = 1'b0;
	assign bitmap[1114] = 1'b1;
	assign bitmap[1115] = 1'b0;
	assign bitmap[1116] = 1'b0;
	assign bitmap[1117] = 1'b1;
	assign bitmap[1118] = 1'b0;
	assign bitmap[1119] = 1'b0;
	assign bitmap[1120] = 1'b0;
	assign bitmap[1121] = 1'b0;
	assign bitmap[1122] = 1'b1;
	assign bitmap[1123] = 1'b1;
	assign bitmap[1124] = 1'b1;
	assign bitmap[1125] = 1'b1;
	assign bitmap[1126] = 1'b0;
	assign bitmap[1127] = 1'b0;
	assign bitmap[1128] = 1'b0;
	assign bitmap[1129] = 1'b0;
	assign bitmap[1130] = 1'b1;
	assign bitmap[1131] = 1'b1;
	assign bitmap[1132] = 1'b1;
	assign bitmap[1133] = 1'b1;
	assign bitmap[1134] = 1'b0;
	assign bitmap[1135] = 1'b0;
	assign bitmap[1136] = 1'b0;
	assign bitmap[1137] = 1'b0;
	assign bitmap[1138] = 1'b0;
	assign bitmap[1139] = 1'b0;
	assign bitmap[1140] = 1'b0;
	assign bitmap[1141] = 1'b0;
	assign bitmap[1142] = 1'b0;
	assign bitmap[1143] = 1'b0;
	assign bitmap[1144] = 1'b0;
	assign bitmap[1145] = 1'b0;
	assign bitmap[1146] = 1'b0;
	assign bitmap[1147] = 1'b0;
	assign bitmap[1148] = 1'b0;
	assign bitmap[1149] = 1'b0;
	assign bitmap[1150] = 1'b0;
	assign bitmap[1151] = 1'b0;
	assign bitmap[1152] = 1'b0;
	assign bitmap[1153] = 1'b0;
	assign bitmap[1154] = 1'b0;
	assign bitmap[1155] = 1'b0;
	assign bitmap[1156] = 1'b0;
	assign bitmap[1157] = 1'b0;
	assign bitmap[1158] = 1'b0;
	assign bitmap[1159] = 1'b0;
	assign bitmap[1160] = 1'b0;
	assign bitmap[1161] = 1'b0;
	assign bitmap[1162] = 1'b0;
	assign bitmap[1163] = 1'b0;
	assign bitmap[1164] = 1'b0;
	assign bitmap[1165] = 1'b0;
	assign bitmap[1166] = 1'b0;
	assign bitmap[1167] = 1'b0;
	assign bitmap[1168] = 1'b0;
	assign bitmap[1169] = 1'b0;
	assign bitmap[1170] = 1'b0;
	assign bitmap[1171] = 1'b0;
	assign bitmap[1172] = 1'b0;
	assign bitmap[1173] = 1'b0;
	assign bitmap[1174] = 1'b0;
	assign bitmap[1175] = 1'b0;
	assign bitmap[1176] = 1'b0;
	assign bitmap[1177] = 1'b0;
	assign bitmap[1178] = 1'b0;
	assign bitmap[1179] = 1'b0;
	assign bitmap[1180] = 1'b0;
	assign bitmap[1181] = 1'b0;
	assign bitmap[1182] = 1'b0;
	assign bitmap[1183] = 1'b0;
	assign bitmap[1184] = 1'b0;
	assign bitmap[1185] = 1'b0;
	assign bitmap[1186] = 1'b0;
	assign bitmap[1187] = 1'b0;
	assign bitmap[1188] = 1'b0;
	assign bitmap[1189] = 1'b0;
	assign bitmap[1190] = 1'b0;
	assign bitmap[1191] = 1'b0;
	assign bitmap[1192] = 1'b0;
	assign bitmap[1193] = 1'b0;
	assign bitmap[1194] = 1'b0;
	assign bitmap[1195] = 1'b0;
	assign bitmap[1196] = 1'b0;
	assign bitmap[1197] = 1'b0;
	assign bitmap[1198] = 1'b0;
	assign bitmap[1199] = 1'b0;
	assign bitmap[1200] = 1'b0;
	assign bitmap[1201] = 1'b0;
	assign bitmap[1202] = 1'b0;
	assign bitmap[1203] = 1'b0;
	assign bitmap[1204] = 1'b0;
	assign bitmap[1205] = 1'b0;
	assign bitmap[1206] = 1'b0;
	assign bitmap[1207] = 1'b0;
	assign bitmap[1208] = 1'b0;
	assign bitmap[1209] = 1'b0;
	assign bitmap[1210] = 1'b0;
	assign bitmap[1211] = 1'b0;
	assign bitmap[1212] = 1'b0;
	assign bitmap[1213] = 1'b0;
	assign bitmap[1214] = 1'b0;
	assign bitmap[1215] = 1'b0;
	assign bitmap[1216] = 1'b0;
	assign bitmap[1217] = 1'b0;
	assign bitmap[1218] = 1'b0;
	assign bitmap[1219] = 1'b0;
	assign bitmap[1220] = 1'b0;
	assign bitmap[1221] = 1'b0;
	assign bitmap[1222] = 1'b0;
	assign bitmap[1223] = 1'b0;
	assign bitmap[1224] = 1'b0;
	assign bitmap[1225] = 1'b0;
	assign bitmap[1226] = 1'b0;
	assign bitmap[1227] = 1'b0;
	assign bitmap[1228] = 1'b0;
	assign bitmap[1229] = 1'b0;
	assign bitmap[1230] = 1'b0;
	assign bitmap[1231] = 1'b0;
	assign bitmap[1232] = 1'b0;
	assign bitmap[1233] = 1'b0;
	assign bitmap[1234] = 1'b0;
	assign bitmap[1235] = 1'b0;
	assign bitmap[1236] = 1'b0;
	assign bitmap[1237] = 1'b0;
	assign bitmap[1238] = 1'b0;
	assign bitmap[1239] = 1'b0;
	assign bitmap[1240] = 1'b0;
	assign bitmap[1241] = 1'b0;
	assign bitmap[1242] = 1'b0;
	assign bitmap[1243] = 1'b0;
	assign bitmap[1244] = 1'b0;
	assign bitmap[1245] = 1'b0;
	assign bitmap[1246] = 1'b0;
	assign bitmap[1247] = 1'b0;
	assign bitmap[1248] = 1'b0;
	assign bitmap[1249] = 1'b0;
	assign bitmap[1250] = 1'b0;
	assign bitmap[1251] = 1'b0;
	assign bitmap[1252] = 1'b0;
	assign bitmap[1253] = 1'b0;
	assign bitmap[1254] = 1'b0;
	assign bitmap[1255] = 1'b0;
	assign bitmap[1256] = 1'b0;
	assign bitmap[1257] = 1'b0;
	assign bitmap[1258] = 1'b0;
	assign bitmap[1259] = 1'b0;
	assign bitmap[1260] = 1'b0;
	assign bitmap[1261] = 1'b0;
	assign bitmap[1262] = 1'b0;
	assign bitmap[1263] = 1'b0;
	assign bitmap[1264] = 1'b0;
	assign bitmap[1265] = 1'b0;
	assign bitmap[1266] = 1'b0;
	assign bitmap[1267] = 1'b0;
	assign bitmap[1268] = 1'b0;
	assign bitmap[1269] = 1'b0;
	assign bitmap[1270] = 1'b0;
	assign bitmap[1271] = 1'b0;
	assign bitmap[1272] = 1'b0;
	assign bitmap[1273] = 1'b0;
	assign bitmap[1274] = 1'b0;
	assign bitmap[1275] = 1'b0;
	assign bitmap[1276] = 1'b0;
	assign bitmap[1277] = 1'b0;
	assign bitmap[1278] = 1'b0;
	assign bitmap[1279] = 1'b0;
	assign bitmap[1280] = 1'b0;
	assign bitmap[1281] = 1'b0;
	assign bitmap[1282] = 1'b0;
	assign bitmap[1283] = 1'b0;
	assign bitmap[1284] = 1'b0;
	assign bitmap[1285] = 1'b0;
	assign bitmap[1286] = 1'b0;
	assign bitmap[1287] = 1'b0;
	assign bitmap[1288] = 1'b0;
	assign bitmap[1289] = 1'b0;
	assign bitmap[1290] = 1'b0;
	assign bitmap[1291] = 1'b0;
	assign bitmap[1292] = 1'b0;
	assign bitmap[1293] = 1'b0;
	assign bitmap[1294] = 1'b0;
	assign bitmap[1295] = 1'b0;
	assign bitmap[1296] = 1'b0;
	assign bitmap[1297] = 1'b0;
	assign bitmap[1298] = 1'b1;
	assign bitmap[1299] = 1'b1;
	assign bitmap[1300] = 1'b1;
	assign bitmap[1301] = 1'b1;
	assign bitmap[1302] = 1'b0;
	assign bitmap[1303] = 1'b0;
	assign bitmap[1304] = 1'b0;
	assign bitmap[1305] = 1'b0;
	assign bitmap[1306] = 1'b0;
	assign bitmap[1307] = 1'b1;
	assign bitmap[1308] = 1'b1;
	assign bitmap[1309] = 1'b0;
	assign bitmap[1310] = 1'b0;
	assign bitmap[1311] = 1'b0;
	assign bitmap[1312] = 1'b0;
	assign bitmap[1313] = 1'b0;
	assign bitmap[1314] = 1'b0;
	assign bitmap[1315] = 1'b0;
	assign bitmap[1316] = 1'b0;
	assign bitmap[1317] = 1'b1;
	assign bitmap[1318] = 1'b0;
	assign bitmap[1319] = 1'b0;
	assign bitmap[1320] = 1'b0;
	assign bitmap[1321] = 1'b0;
	assign bitmap[1322] = 1'b1;
	assign bitmap[1323] = 1'b0;
	assign bitmap[1324] = 1'b0;
	assign bitmap[1325] = 1'b1;
	assign bitmap[1326] = 1'b0;
	assign bitmap[1327] = 1'b0;
	assign bitmap[1328] = 1'b0;
	assign bitmap[1329] = 1'b0;
	assign bitmap[1330] = 1'b0;
	assign bitmap[1331] = 1'b0;
	assign bitmap[1332] = 1'b0;
	assign bitmap[1333] = 1'b1;
	assign bitmap[1334] = 1'b0;
	assign bitmap[1335] = 1'b0;
	assign bitmap[1336] = 1'b0;
	assign bitmap[1337] = 1'b0;
	assign bitmap[1338] = 1'b0;
	assign bitmap[1339] = 1'b0;
	assign bitmap[1340] = 1'b0;
	assign bitmap[1341] = 1'b1;
	assign bitmap[1342] = 1'b0;
	assign bitmap[1343] = 1'b0;
	assign bitmap[1344] = 1'b0;
	assign bitmap[1345] = 1'b0;
	assign bitmap[1346] = 1'b1;
	assign bitmap[1347] = 1'b1;
	assign bitmap[1348] = 1'b1;
	assign bitmap[1349] = 1'b1;
	assign bitmap[1350] = 1'b0;
	assign bitmap[1351] = 1'b0;
	assign bitmap[1352] = 1'b0;
	assign bitmap[1353] = 1'b0;
	assign bitmap[1354] = 1'b0;
	assign bitmap[1355] = 1'b0;
	assign bitmap[1356] = 1'b1;
	assign bitmap[1357] = 1'b0;
	assign bitmap[1358] = 1'b0;
	assign bitmap[1359] = 1'b0;
	assign bitmap[1360] = 1'b0;
	assign bitmap[1361] = 1'b0;
	assign bitmap[1362] = 1'b0;
	assign bitmap[1363] = 1'b0;
	assign bitmap[1364] = 1'b0;
	assign bitmap[1365] = 1'b1;
	assign bitmap[1366] = 1'b0;
	assign bitmap[1367] = 1'b0;
	assign bitmap[1368] = 1'b0;
	assign bitmap[1369] = 1'b0;
	assign bitmap[1370] = 1'b0;
	assign bitmap[1371] = 1'b1;
	assign bitmap[1372] = 1'b0;
	assign bitmap[1373] = 1'b0;
	assign bitmap[1374] = 1'b0;
	assign bitmap[1375] = 1'b0;
	assign bitmap[1376] = 1'b0;
	assign bitmap[1377] = 1'b0;
	assign bitmap[1378] = 1'b1;
	assign bitmap[1379] = 1'b1;
	assign bitmap[1380] = 1'b1;
	assign bitmap[1381] = 1'b1;
	assign bitmap[1382] = 1'b0;
	assign bitmap[1383] = 1'b0;
	assign bitmap[1384] = 1'b0;
	assign bitmap[1385] = 1'b0;
	assign bitmap[1386] = 1'b1;
	assign bitmap[1387] = 1'b1;
	assign bitmap[1388] = 1'b1;
	assign bitmap[1389] = 1'b1;
	assign bitmap[1390] = 1'b0;
	assign bitmap[1391] = 1'b0;
	assign bitmap[1392] = 1'b0;
	assign bitmap[1393] = 1'b0;
	assign bitmap[1394] = 1'b0;
	assign bitmap[1395] = 1'b0;
	assign bitmap[1396] = 1'b0;
	assign bitmap[1397] = 1'b0;
	assign bitmap[1398] = 1'b0;
	assign bitmap[1399] = 1'b0;
	assign bitmap[1400] = 1'b0;
	assign bitmap[1401] = 1'b0;
	assign bitmap[1402] = 1'b0;
	assign bitmap[1403] = 1'b0;
	assign bitmap[1404] = 1'b0;
	assign bitmap[1405] = 1'b0;
	assign bitmap[1406] = 1'b0;
	assign bitmap[1407] = 1'b0;
	assign bitmap[1408] = 1'b0;
	assign bitmap[1409] = 1'b0;
	assign bitmap[1410] = 1'b0;
	assign bitmap[1411] = 1'b0;
	assign bitmap[1412] = 1'b0;
	assign bitmap[1413] = 1'b0;
	assign bitmap[1414] = 1'b0;
	assign bitmap[1415] = 1'b0;
	assign bitmap[1416] = 1'b0;
	assign bitmap[1417] = 1'b0;
	assign bitmap[1418] = 1'b0;
	assign bitmap[1419] = 1'b0;
	assign bitmap[1420] = 1'b0;
	assign bitmap[1421] = 1'b0;
	assign bitmap[1422] = 1'b0;
	assign bitmap[1423] = 1'b0;
	assign bitmap[1424] = 1'b0;
	assign bitmap[1425] = 1'b0;
	assign bitmap[1426] = 1'b0;
	assign bitmap[1427] = 1'b0;
	assign bitmap[1428] = 1'b0;
	assign bitmap[1429] = 1'b0;
	assign bitmap[1430] = 1'b0;
	assign bitmap[1431] = 1'b0;
	assign bitmap[1432] = 1'b0;
	assign bitmap[1433] = 1'b0;
	assign bitmap[1434] = 1'b0;
	assign bitmap[1435] = 1'b0;
	assign bitmap[1436] = 1'b0;
	assign bitmap[1437] = 1'b0;
	assign bitmap[1438] = 1'b0;
	assign bitmap[1439] = 1'b0;
	assign bitmap[1440] = 1'b0;
	assign bitmap[1441] = 1'b0;
	assign bitmap[1442] = 1'b0;
	assign bitmap[1443] = 1'b0;
	assign bitmap[1444] = 1'b0;
	assign bitmap[1445] = 1'b0;
	assign bitmap[1446] = 1'b0;
	assign bitmap[1447] = 1'b0;
	assign bitmap[1448] = 1'b0;
	assign bitmap[1449] = 1'b0;
	assign bitmap[1450] = 1'b0;
	assign bitmap[1451] = 1'b0;
	assign bitmap[1452] = 1'b0;
	assign bitmap[1453] = 1'b0;
	assign bitmap[1454] = 1'b0;
	assign bitmap[1455] = 1'b0;
	assign bitmap[1456] = 1'b0;
	assign bitmap[1457] = 1'b0;
	assign bitmap[1458] = 1'b0;
	assign bitmap[1459] = 1'b0;
	assign bitmap[1460] = 1'b0;
	assign bitmap[1461] = 1'b0;
	assign bitmap[1462] = 1'b0;
	assign bitmap[1463] = 1'b0;
	assign bitmap[1464] = 1'b0;
	assign bitmap[1465] = 1'b0;
	assign bitmap[1466] = 1'b0;
	assign bitmap[1467] = 1'b0;
	assign bitmap[1468] = 1'b0;
	assign bitmap[1469] = 1'b0;
	assign bitmap[1470] = 1'b0;
	assign bitmap[1471] = 1'b0;
	assign bitmap[1472] = 1'b0;
	assign bitmap[1473] = 1'b0;
	assign bitmap[1474] = 1'b0;
	assign bitmap[1475] = 1'b0;
	assign bitmap[1476] = 1'b0;
	assign bitmap[1477] = 1'b0;
	assign bitmap[1478] = 1'b0;
	assign bitmap[1479] = 1'b0;
	assign bitmap[1480] = 1'b0;
	assign bitmap[1481] = 1'b0;
	assign bitmap[1482] = 1'b0;
	assign bitmap[1483] = 1'b0;
	assign bitmap[1484] = 1'b0;
	assign bitmap[1485] = 1'b0;
	assign bitmap[1486] = 1'b0;
	assign bitmap[1487] = 1'b0;
	assign bitmap[1488] = 1'b0;
	assign bitmap[1489] = 1'b0;
	assign bitmap[1490] = 1'b0;
	assign bitmap[1491] = 1'b0;
	assign bitmap[1492] = 1'b0;
	assign bitmap[1493] = 1'b0;
	assign bitmap[1494] = 1'b0;
	assign bitmap[1495] = 1'b0;
	assign bitmap[1496] = 1'b0;
	assign bitmap[1497] = 1'b0;
	assign bitmap[1498] = 1'b0;
	assign bitmap[1499] = 1'b0;
	assign bitmap[1500] = 1'b0;
	assign bitmap[1501] = 1'b0;
	assign bitmap[1502] = 1'b0;
	assign bitmap[1503] = 1'b0;
	assign bitmap[1504] = 1'b0;
	assign bitmap[1505] = 1'b0;
	assign bitmap[1506] = 1'b0;
	assign bitmap[1507] = 1'b0;
	assign bitmap[1508] = 1'b0;
	assign bitmap[1509] = 1'b0;
	assign bitmap[1510] = 1'b0;
	assign bitmap[1511] = 1'b0;
	assign bitmap[1512] = 1'b0;
	assign bitmap[1513] = 1'b0;
	assign bitmap[1514] = 1'b0;
	assign bitmap[1515] = 1'b0;
	assign bitmap[1516] = 1'b0;
	assign bitmap[1517] = 1'b0;
	assign bitmap[1518] = 1'b0;
	assign bitmap[1519] = 1'b0;
	assign bitmap[1520] = 1'b0;
	assign bitmap[1521] = 1'b0;
	assign bitmap[1522] = 1'b0;
	assign bitmap[1523] = 1'b0;
	assign bitmap[1524] = 1'b0;
	assign bitmap[1525] = 1'b0;
	assign bitmap[1526] = 1'b0;
	assign bitmap[1527] = 1'b0;
	assign bitmap[1528] = 1'b0;
	assign bitmap[1529] = 1'b0;
	assign bitmap[1530] = 1'b0;
	assign bitmap[1531] = 1'b0;
	assign bitmap[1532] = 1'b0;
	assign bitmap[1533] = 1'b0;
	assign bitmap[1534] = 1'b0;
	assign bitmap[1535] = 1'b0;
	assign bitmap[1536] = 1'b0;
	assign bitmap[1537] = 1'b0;
	assign bitmap[1538] = 1'b0;
	assign bitmap[1539] = 1'b0;
	assign bitmap[1540] = 1'b0;
	assign bitmap[1541] = 1'b0;
	assign bitmap[1542] = 1'b0;
	assign bitmap[1543] = 1'b0;
	assign bitmap[1544] = 1'b0;
	assign bitmap[1545] = 1'b0;
	assign bitmap[1546] = 1'b0;
	assign bitmap[1547] = 1'b0;
	assign bitmap[1548] = 1'b0;
	assign bitmap[1549] = 1'b0;
	assign bitmap[1550] = 1'b0;
	assign bitmap[1551] = 1'b0;
	assign bitmap[1552] = 1'b0;
	assign bitmap[1553] = 1'b0;
	assign bitmap[1554] = 1'b1;
	assign bitmap[1555] = 1'b1;
	assign bitmap[1556] = 1'b1;
	assign bitmap[1557] = 1'b1;
	assign bitmap[1558] = 1'b0;
	assign bitmap[1559] = 1'b0;
	assign bitmap[1560] = 1'b0;
	assign bitmap[1561] = 1'b0;
	assign bitmap[1562] = 1'b0;
	assign bitmap[1563] = 1'b0;
	assign bitmap[1564] = 1'b1;
	assign bitmap[1565] = 1'b1;
	assign bitmap[1566] = 1'b0;
	assign bitmap[1567] = 1'b0;
	assign bitmap[1568] = 1'b0;
	assign bitmap[1569] = 1'b0;
	assign bitmap[1570] = 1'b1;
	assign bitmap[1571] = 1'b0;
	assign bitmap[1572] = 1'b0;
	assign bitmap[1573] = 1'b0;
	assign bitmap[1574] = 1'b0;
	assign bitmap[1575] = 1'b0;
	assign bitmap[1576] = 1'b0;
	assign bitmap[1577] = 1'b0;
	assign bitmap[1578] = 1'b0;
	assign bitmap[1579] = 1'b1;
	assign bitmap[1580] = 1'b0;
	assign bitmap[1581] = 1'b1;
	assign bitmap[1582] = 1'b0;
	assign bitmap[1583] = 1'b0;
	assign bitmap[1584] = 1'b0;
	assign bitmap[1585] = 1'b0;
	assign bitmap[1586] = 1'b1;
	assign bitmap[1587] = 1'b0;
	assign bitmap[1588] = 1'b0;
	assign bitmap[1589] = 1'b0;
	assign bitmap[1590] = 1'b0;
	assign bitmap[1591] = 1'b0;
	assign bitmap[1592] = 1'b0;
	assign bitmap[1593] = 1'b0;
	assign bitmap[1594] = 1'b1;
	assign bitmap[1595] = 1'b0;
	assign bitmap[1596] = 1'b0;
	assign bitmap[1597] = 1'b1;
	assign bitmap[1598] = 1'b0;
	assign bitmap[1599] = 1'b0;
	assign bitmap[1600] = 1'b0;
	assign bitmap[1601] = 1'b0;
	assign bitmap[1602] = 1'b1;
	assign bitmap[1603] = 1'b1;
	assign bitmap[1604] = 1'b1;
	assign bitmap[1605] = 1'b1;
	assign bitmap[1606] = 1'b0;
	assign bitmap[1607] = 1'b0;
	assign bitmap[1608] = 1'b0;
	assign bitmap[1609] = 1'b0;
	assign bitmap[1610] = 1'b1;
	assign bitmap[1611] = 1'b1;
	assign bitmap[1612] = 1'b1;
	assign bitmap[1613] = 1'b1;
	assign bitmap[1614] = 1'b1;
	assign bitmap[1615] = 1'b0;
	assign bitmap[1616] = 1'b0;
	assign bitmap[1617] = 1'b0;
	assign bitmap[1618] = 1'b1;
	assign bitmap[1619] = 1'b0;
	assign bitmap[1620] = 1'b0;
	assign bitmap[1621] = 1'b1;
	assign bitmap[1622] = 1'b0;
	assign bitmap[1623] = 1'b0;
	assign bitmap[1624] = 1'b0;
	assign bitmap[1625] = 1'b0;
	assign bitmap[1626] = 1'b0;
	assign bitmap[1627] = 1'b0;
	assign bitmap[1628] = 1'b0;
	assign bitmap[1629] = 1'b1;
	assign bitmap[1630] = 1'b0;
	assign bitmap[1631] = 1'b0;
	assign bitmap[1632] = 1'b0;
	assign bitmap[1633] = 1'b0;
	assign bitmap[1634] = 1'b1;
	assign bitmap[1635] = 1'b1;
	assign bitmap[1636] = 1'b1;
	assign bitmap[1637] = 1'b1;
	assign bitmap[1638] = 1'b0;
	assign bitmap[1639] = 1'b0;
	assign bitmap[1640] = 1'b0;
	assign bitmap[1641] = 1'b0;
	assign bitmap[1642] = 1'b0;
	assign bitmap[1643] = 1'b0;
	assign bitmap[1644] = 1'b0;
	assign bitmap[1645] = 1'b1;
	assign bitmap[1646] = 1'b0;
	assign bitmap[1647] = 1'b0;
	assign bitmap[1648] = 1'b0;
	assign bitmap[1649] = 1'b0;
	assign bitmap[1650] = 1'b0;
	assign bitmap[1651] = 1'b0;
	assign bitmap[1652] = 1'b0;
	assign bitmap[1653] = 1'b0;
	assign bitmap[1654] = 1'b0;
	assign bitmap[1655] = 1'b0;
	assign bitmap[1656] = 1'b0;
	assign bitmap[1657] = 1'b0;
	assign bitmap[1658] = 1'b0;
	assign bitmap[1659] = 1'b0;
	assign bitmap[1660] = 1'b0;
	assign bitmap[1661] = 1'b0;
	assign bitmap[1662] = 1'b0;
	assign bitmap[1663] = 1'b0;
	assign bitmap[1664] = 1'b0;
	assign bitmap[1665] = 1'b0;
	assign bitmap[1666] = 1'b0;
	assign bitmap[1667] = 1'b0;
	assign bitmap[1668] = 1'b0;
	assign bitmap[1669] = 1'b0;
	assign bitmap[1670] = 1'b0;
	assign bitmap[1671] = 1'b0;
	assign bitmap[1672] = 1'b0;
	assign bitmap[1673] = 1'b0;
	assign bitmap[1674] = 1'b0;
	assign bitmap[1675] = 1'b0;
	assign bitmap[1676] = 1'b0;
	assign bitmap[1677] = 1'b0;
	assign bitmap[1678] = 1'b0;
	assign bitmap[1679] = 1'b0;
	assign bitmap[1680] = 1'b0;
	assign bitmap[1681] = 1'b0;
	assign bitmap[1682] = 1'b0;
	assign bitmap[1683] = 1'b0;
	assign bitmap[1684] = 1'b0;
	assign bitmap[1685] = 1'b0;
	assign bitmap[1686] = 1'b0;
	assign bitmap[1687] = 1'b0;
	assign bitmap[1688] = 1'b0;
	assign bitmap[1689] = 1'b0;
	assign bitmap[1690] = 1'b0;
	assign bitmap[1691] = 1'b0;
	assign bitmap[1692] = 1'b0;
	assign bitmap[1693] = 1'b0;
	assign bitmap[1694] = 1'b0;
	assign bitmap[1695] = 1'b0;
	assign bitmap[1696] = 1'b0;
	assign bitmap[1697] = 1'b0;
	assign bitmap[1698] = 1'b0;
	assign bitmap[1699] = 1'b0;
	assign bitmap[1700] = 1'b0;
	assign bitmap[1701] = 1'b0;
	assign bitmap[1702] = 1'b0;
	assign bitmap[1703] = 1'b0;
	assign bitmap[1704] = 1'b0;
	assign bitmap[1705] = 1'b0;
	assign bitmap[1706] = 1'b0;
	assign bitmap[1707] = 1'b0;
	assign bitmap[1708] = 1'b0;
	assign bitmap[1709] = 1'b0;
	assign bitmap[1710] = 1'b0;
	assign bitmap[1711] = 1'b0;
	assign bitmap[1712] = 1'b0;
	assign bitmap[1713] = 1'b0;
	assign bitmap[1714] = 1'b0;
	assign bitmap[1715] = 1'b0;
	assign bitmap[1716] = 1'b0;
	assign bitmap[1717] = 1'b0;
	assign bitmap[1718] = 1'b0;
	assign bitmap[1719] = 1'b0;
	assign bitmap[1720] = 1'b0;
	assign bitmap[1721] = 1'b0;
	assign bitmap[1722] = 1'b0;
	assign bitmap[1723] = 1'b0;
	assign bitmap[1724] = 1'b0;
	assign bitmap[1725] = 1'b0;
	assign bitmap[1726] = 1'b0;
	assign bitmap[1727] = 1'b0;
	assign bitmap[1728] = 1'b0;
	assign bitmap[1729] = 1'b0;
	assign bitmap[1730] = 1'b0;
	assign bitmap[1731] = 1'b0;
	assign bitmap[1732] = 1'b0;
	assign bitmap[1733] = 1'b0;
	assign bitmap[1734] = 1'b0;
	assign bitmap[1735] = 1'b0;
	assign bitmap[1736] = 1'b0;
	assign bitmap[1737] = 1'b0;
	assign bitmap[1738] = 1'b0;
	assign bitmap[1739] = 1'b0;
	assign bitmap[1740] = 1'b0;
	assign bitmap[1741] = 1'b0;
	assign bitmap[1742] = 1'b0;
	assign bitmap[1743] = 1'b0;
	assign bitmap[1744] = 1'b0;
	assign bitmap[1745] = 1'b0;
	assign bitmap[1746] = 1'b0;
	assign bitmap[1747] = 1'b0;
	assign bitmap[1748] = 1'b0;
	assign bitmap[1749] = 1'b0;
	assign bitmap[1750] = 1'b0;
	assign bitmap[1751] = 1'b0;
	assign bitmap[1752] = 1'b0;
	assign bitmap[1753] = 1'b0;
	assign bitmap[1754] = 1'b0;
	assign bitmap[1755] = 1'b0;
	assign bitmap[1756] = 1'b0;
	assign bitmap[1757] = 1'b0;
	assign bitmap[1758] = 1'b0;
	assign bitmap[1759] = 1'b0;
	assign bitmap[1760] = 1'b0;
	assign bitmap[1761] = 1'b0;
	assign bitmap[1762] = 1'b0;
	assign bitmap[1763] = 1'b0;
	assign bitmap[1764] = 1'b0;
	assign bitmap[1765] = 1'b0;
	assign bitmap[1766] = 1'b0;
	assign bitmap[1767] = 1'b0;
	assign bitmap[1768] = 1'b0;
	assign bitmap[1769] = 1'b0;
	assign bitmap[1770] = 1'b0;
	assign bitmap[1771] = 1'b0;
	assign bitmap[1772] = 1'b0;
	assign bitmap[1773] = 1'b0;
	assign bitmap[1774] = 1'b0;
	assign bitmap[1775] = 1'b0;
	assign bitmap[1776] = 1'b0;
	assign bitmap[1777] = 1'b0;
	assign bitmap[1778] = 1'b0;
	assign bitmap[1779] = 1'b0;
	assign bitmap[1780] = 1'b0;
	assign bitmap[1781] = 1'b0;
	assign bitmap[1782] = 1'b0;
	assign bitmap[1783] = 1'b0;
	assign bitmap[1784] = 1'b0;
	assign bitmap[1785] = 1'b0;
	assign bitmap[1786] = 1'b0;
	assign bitmap[1787] = 1'b0;
	assign bitmap[1788] = 1'b0;
	assign bitmap[1789] = 1'b0;
	assign bitmap[1790] = 1'b0;
	assign bitmap[1791] = 1'b0;
	assign bitmap[1792] = 1'b0;
	assign bitmap[1793] = 1'b0;
	assign bitmap[1794] = 1'b0;
	assign bitmap[1795] = 1'b0;
	assign bitmap[1796] = 1'b0;
	assign bitmap[1797] = 1'b0;
	assign bitmap[1798] = 1'b0;
	assign bitmap[1799] = 1'b0;
	assign bitmap[1800] = 1'b0;
	assign bitmap[1801] = 1'b0;
	assign bitmap[1802] = 1'b0;
	assign bitmap[1803] = 1'b0;
	assign bitmap[1804] = 1'b0;
	assign bitmap[1805] = 1'b0;
	assign bitmap[1806] = 1'b0;
	assign bitmap[1807] = 1'b0;
	assign bitmap[1808] = 1'b0;
	assign bitmap[1809] = 1'b0;
	assign bitmap[1810] = 1'b0;
	assign bitmap[1811] = 1'b0;
	assign bitmap[1812] = 1'b1;
	assign bitmap[1813] = 1'b0;
	assign bitmap[1814] = 1'b0;
	assign bitmap[1815] = 1'b0;
	assign bitmap[1816] = 1'b0;
	assign bitmap[1817] = 1'b0;
	assign bitmap[1818] = 1'b0;
	assign bitmap[1819] = 1'b1;
	assign bitmap[1820] = 1'b1;
	assign bitmap[1821] = 1'b0;
	assign bitmap[1822] = 1'b0;
	assign bitmap[1823] = 1'b0;
	assign bitmap[1824] = 1'b0;
	assign bitmap[1825] = 1'b0;
	assign bitmap[1826] = 1'b0;
	assign bitmap[1827] = 1'b1;
	assign bitmap[1828] = 1'b1;
	assign bitmap[1829] = 1'b0;
	assign bitmap[1830] = 1'b0;
	assign bitmap[1831] = 1'b0;
	assign bitmap[1832] = 1'b0;
	assign bitmap[1833] = 1'b0;
	assign bitmap[1834] = 1'b1;
	assign bitmap[1835] = 1'b0;
	assign bitmap[1836] = 1'b0;
	assign bitmap[1837] = 1'b1;
	assign bitmap[1838] = 1'b0;
	assign bitmap[1839] = 1'b0;
	assign bitmap[1840] = 1'b0;
	assign bitmap[1841] = 1'b0;
	assign bitmap[1842] = 1'b1;
	assign bitmap[1843] = 1'b0;
	assign bitmap[1844] = 1'b1;
	assign bitmap[1845] = 1'b0;
	assign bitmap[1846] = 1'b0;
	assign bitmap[1847] = 1'b0;
	assign bitmap[1848] = 1'b0;
	assign bitmap[1849] = 1'b0;
	assign bitmap[1850] = 1'b0;
	assign bitmap[1851] = 1'b0;
	assign bitmap[1852] = 1'b0;
	assign bitmap[1853] = 1'b1;
	assign bitmap[1854] = 1'b0;
	assign bitmap[1855] = 1'b0;
	assign bitmap[1856] = 1'b0;
	assign bitmap[1857] = 1'b0;
	assign bitmap[1858] = 1'b0;
	assign bitmap[1859] = 1'b0;
	assign bitmap[1860] = 1'b1;
	assign bitmap[1861] = 1'b0;
	assign bitmap[1862] = 1'b0;
	assign bitmap[1863] = 1'b0;
	assign bitmap[1864] = 1'b0;
	assign bitmap[1865] = 1'b0;
	assign bitmap[1866] = 1'b0;
	assign bitmap[1867] = 1'b0;
	assign bitmap[1868] = 1'b1;
	assign bitmap[1869] = 1'b0;
	assign bitmap[1870] = 1'b0;
	assign bitmap[1871] = 1'b0;
	assign bitmap[1872] = 1'b0;
	assign bitmap[1873] = 1'b0;
	assign bitmap[1874] = 1'b0;
	assign bitmap[1875] = 1'b0;
	assign bitmap[1876] = 1'b1;
	assign bitmap[1877] = 1'b0;
	assign bitmap[1878] = 1'b0;
	assign bitmap[1879] = 1'b0;
	assign bitmap[1880] = 1'b0;
	assign bitmap[1881] = 1'b0;
	assign bitmap[1882] = 1'b0;
	assign bitmap[1883] = 1'b1;
	assign bitmap[1884] = 1'b0;
	assign bitmap[1885] = 1'b0;
	assign bitmap[1886] = 1'b0;
	assign bitmap[1887] = 1'b0;
	assign bitmap[1888] = 1'b0;
	assign bitmap[1889] = 1'b0;
	assign bitmap[1890] = 1'b1;
	assign bitmap[1891] = 1'b1;
	assign bitmap[1892] = 1'b1;
	assign bitmap[1893] = 1'b1;
	assign bitmap[1894] = 1'b0;
	assign bitmap[1895] = 1'b0;
	assign bitmap[1896] = 1'b0;
	assign bitmap[1897] = 1'b0;
	assign bitmap[1898] = 1'b1;
	assign bitmap[1899] = 1'b1;
	assign bitmap[1900] = 1'b1;
	assign bitmap[1901] = 1'b1;
	assign bitmap[1902] = 1'b0;
	assign bitmap[1903] = 1'b0;
	assign bitmap[1904] = 1'b0;
	assign bitmap[1905] = 1'b0;
	assign bitmap[1906] = 1'b0;
	assign bitmap[1907] = 1'b0;
	assign bitmap[1908] = 1'b0;
	assign bitmap[1909] = 1'b0;
	assign bitmap[1910] = 1'b0;
	assign bitmap[1911] = 1'b0;
	assign bitmap[1912] = 1'b0;
	assign bitmap[1913] = 1'b0;
	assign bitmap[1914] = 1'b0;
	assign bitmap[1915] = 1'b0;
	assign bitmap[1916] = 1'b0;
	assign bitmap[1917] = 1'b0;
	assign bitmap[1918] = 1'b0;
	assign bitmap[1919] = 1'b0;
	assign bitmap[1920] = 1'b0;
	assign bitmap[1921] = 1'b0;
	assign bitmap[1922] = 1'b0;
	assign bitmap[1923] = 1'b0;
	assign bitmap[1924] = 1'b0;
	assign bitmap[1925] = 1'b0;
	assign bitmap[1926] = 1'b0;
	assign bitmap[1927] = 1'b0;
	assign bitmap[1928] = 1'b0;
	assign bitmap[1929] = 1'b0;
	assign bitmap[1930] = 1'b0;
	assign bitmap[1931] = 1'b0;
	assign bitmap[1932] = 1'b0;
	assign bitmap[1933] = 1'b0;
	assign bitmap[1934] = 1'b0;
	assign bitmap[1935] = 1'b0;
	assign bitmap[1936] = 1'b0;
	assign bitmap[1937] = 1'b0;
	assign bitmap[1938] = 1'b1;
	assign bitmap[1939] = 1'b1;
	assign bitmap[1940] = 1'b1;
	assign bitmap[1941] = 1'b1;
	assign bitmap[1942] = 1'b0;
	assign bitmap[1943] = 1'b0;
	assign bitmap[1944] = 1'b0;
	assign bitmap[1945] = 1'b0;
	assign bitmap[1946] = 1'b0;
	assign bitmap[1947] = 1'b0;
	assign bitmap[1948] = 1'b0;
	assign bitmap[1949] = 1'b0;
	assign bitmap[1950] = 1'b0;
	assign bitmap[1951] = 1'b0;
	assign bitmap[1952] = 1'b0;
	assign bitmap[1953] = 1'b0;
	assign bitmap[1954] = 1'b1;
	assign bitmap[1955] = 1'b0;
	assign bitmap[1956] = 1'b0;
	assign bitmap[1957] = 1'b1;
	assign bitmap[1958] = 1'b0;
	assign bitmap[1959] = 1'b0;
	assign bitmap[1960] = 1'b0;
	assign bitmap[1961] = 1'b0;
	assign bitmap[1962] = 1'b0;
	assign bitmap[1963] = 1'b0;
	assign bitmap[1964] = 1'b0;
	assign bitmap[1965] = 1'b0;
	assign bitmap[1966] = 1'b0;
	assign bitmap[1967] = 1'b0;
	assign bitmap[1968] = 1'b0;
	assign bitmap[1969] = 1'b0;
	assign bitmap[1970] = 1'b1;
	assign bitmap[1971] = 1'b0;
	assign bitmap[1972] = 1'b0;
	assign bitmap[1973] = 1'b1;
	assign bitmap[1974] = 1'b0;
	assign bitmap[1975] = 1'b0;
	assign bitmap[1976] = 1'b0;
	assign bitmap[1977] = 1'b0;
	assign bitmap[1978] = 1'b0;
	assign bitmap[1979] = 1'b0;
	assign bitmap[1980] = 1'b0;
	assign bitmap[1981] = 1'b0;
	assign bitmap[1982] = 1'b0;
	assign bitmap[1983] = 1'b0;
	assign bitmap[1984] = 1'b0;
	assign bitmap[1985] = 1'b0;
	assign bitmap[1986] = 1'b1;
	assign bitmap[1987] = 1'b1;
	assign bitmap[1988] = 1'b1;
	assign bitmap[1989] = 1'b1;
	assign bitmap[1990] = 1'b0;
	assign bitmap[1991] = 1'b0;
	assign bitmap[1992] = 1'b0;
	assign bitmap[1993] = 1'b0;
	assign bitmap[1994] = 1'b0;
	assign bitmap[1995] = 1'b0;
	assign bitmap[1996] = 1'b0;
	assign bitmap[1997] = 1'b0;
	assign bitmap[1998] = 1'b0;
	assign bitmap[1999] = 1'b0;
	assign bitmap[2000] = 1'b0;
	assign bitmap[2001] = 1'b0;
	assign bitmap[2002] = 1'b1;
	assign bitmap[2003] = 1'b0;
	assign bitmap[2004] = 1'b0;
	assign bitmap[2005] = 1'b1;
	assign bitmap[2006] = 1'b0;
	assign bitmap[2007] = 1'b0;
	assign bitmap[2008] = 1'b0;
	assign bitmap[2009] = 1'b0;
	assign bitmap[2010] = 1'b0;
	assign bitmap[2011] = 1'b0;
	assign bitmap[2012] = 1'b0;
	assign bitmap[2013] = 1'b0;
	assign bitmap[2014] = 1'b0;
	assign bitmap[2015] = 1'b0;
	assign bitmap[2016] = 1'b0;
	assign bitmap[2017] = 1'b0;
	assign bitmap[2018] = 1'b1;
	assign bitmap[2019] = 1'b1;
	assign bitmap[2020] = 1'b1;
	assign bitmap[2021] = 1'b1;
	assign bitmap[2022] = 1'b0;
	assign bitmap[2023] = 1'b0;
	assign bitmap[2024] = 1'b0;
	assign bitmap[2025] = 1'b0;
	assign bitmap[2026] = 1'b0;
	assign bitmap[2027] = 1'b0;
	assign bitmap[2028] = 1'b0;
	assign bitmap[2029] = 1'b0;
	assign bitmap[2030] = 1'b0;
	assign bitmap[2031] = 1'b0;
	assign bitmap[2032] = 1'b0;
	assign bitmap[2033] = 1'b0;
	assign bitmap[2034] = 1'b0;
	assign bitmap[2035] = 1'b0;
	assign bitmap[2036] = 1'b0;
	assign bitmap[2037] = 1'b0;
	assign bitmap[2038] = 1'b0;
	assign bitmap[2039] = 1'b0;
	assign bitmap[2040] = 1'b0;
	assign bitmap[2041] = 1'b0;
	assign bitmap[2042] = 1'b0;
	assign bitmap[2043] = 1'b0;
	assign bitmap[2044] = 1'b0;
	assign bitmap[2045] = 1'b0;
	assign bitmap[2046] = 1'b0;
	assign bitmap[2047] = 1'b0;
	assign bitmap[2048] = 1'b0;
	assign bitmap[2049] = 1'b0;
	assign bitmap[2050] = 1'b0;
	assign bitmap[2051] = 1'b0;
	assign bitmap[2052] = 1'b0;
	assign bitmap[2053] = 1'b0;
	assign bitmap[2054] = 1'b0;
	assign bitmap[2055] = 1'b0;
	assign bitmap[2056] = 1'b0;
	assign bitmap[2057] = 1'b0;
	assign bitmap[2058] = 1'b0;
	assign bitmap[2059] = 1'b0;
	assign bitmap[2060] = 1'b0;
	assign bitmap[2061] = 1'b0;
	assign bitmap[2062] = 1'b0;
	assign bitmap[2063] = 1'b0;
	assign bitmap[2064] = 1'b0;
	assign bitmap[2065] = 1'b0;
	assign bitmap[2066] = 1'b0;
	assign bitmap[2067] = 1'b1;
	assign bitmap[2068] = 1'b1;
	assign bitmap[2069] = 1'b0;
	assign bitmap[2070] = 1'b0;
	assign bitmap[2071] = 1'b0;
	assign bitmap[2072] = 1'b0;
	assign bitmap[2073] = 1'b0;
	assign bitmap[2074] = 1'b1;
	assign bitmap[2075] = 1'b1;
	assign bitmap[2076] = 1'b1;
	assign bitmap[2077] = 1'b1;
	assign bitmap[2078] = 1'b0;
	assign bitmap[2079] = 1'b0;
	assign bitmap[2080] = 1'b0;
	assign bitmap[2081] = 1'b0;
	assign bitmap[2082] = 1'b1;
	assign bitmap[2083] = 1'b0;
	assign bitmap[2084] = 1'b0;
	assign bitmap[2085] = 1'b1;
	assign bitmap[2086] = 1'b0;
	assign bitmap[2087] = 1'b0;
	assign bitmap[2088] = 1'b0;
	assign bitmap[2089] = 1'b0;
	assign bitmap[2090] = 1'b1;
	assign bitmap[2091] = 1'b0;
	assign bitmap[2092] = 1'b0;
	assign bitmap[2093] = 1'b0;
	assign bitmap[2094] = 1'b0;
	assign bitmap[2095] = 1'b0;
	assign bitmap[2096] = 1'b0;
	assign bitmap[2097] = 1'b0;
	assign bitmap[2098] = 1'b0;
	assign bitmap[2099] = 1'b0;
	assign bitmap[2100] = 1'b0;
	assign bitmap[2101] = 1'b1;
	assign bitmap[2102] = 1'b0;
	assign bitmap[2103] = 1'b0;
	assign bitmap[2104] = 1'b0;
	assign bitmap[2105] = 1'b0;
	assign bitmap[2106] = 1'b1;
	assign bitmap[2107] = 1'b0;
	assign bitmap[2108] = 1'b0;
	assign bitmap[2109] = 1'b0;
	assign bitmap[2110] = 1'b0;
	assign bitmap[2111] = 1'b0;
	assign bitmap[2112] = 1'b0;
	assign bitmap[2113] = 1'b0;
	assign bitmap[2114] = 1'b0;
	assign bitmap[2115] = 1'b0;
	assign bitmap[2116] = 1'b1;
	assign bitmap[2117] = 1'b0;
	assign bitmap[2118] = 1'b0;
	assign bitmap[2119] = 1'b0;
	assign bitmap[2120] = 1'b0;
	assign bitmap[2121] = 1'b0;
	assign bitmap[2122] = 1'b1;
	assign bitmap[2123] = 1'b1;
	assign bitmap[2124] = 1'b1;
	assign bitmap[2125] = 1'b1;
	assign bitmap[2126] = 1'b0;
	assign bitmap[2127] = 1'b0;
	assign bitmap[2128] = 1'b0;
	assign bitmap[2129] = 1'b0;
	assign bitmap[2130] = 1'b0;
	assign bitmap[2131] = 1'b1;
	assign bitmap[2132] = 1'b0;
	assign bitmap[2133] = 1'b0;
	assign bitmap[2134] = 1'b0;
	assign bitmap[2135] = 1'b0;
	assign bitmap[2136] = 1'b0;
	assign bitmap[2137] = 1'b0;
	assign bitmap[2138] = 1'b0;
	assign bitmap[2139] = 1'b0;
	assign bitmap[2140] = 1'b0;
	assign bitmap[2141] = 1'b1;
	assign bitmap[2142] = 1'b0;
	assign bitmap[2143] = 1'b0;
	assign bitmap[2144] = 1'b0;
	assign bitmap[2145] = 1'b0;
	assign bitmap[2146] = 1'b1;
	assign bitmap[2147] = 1'b1;
	assign bitmap[2148] = 1'b1;
	assign bitmap[2149] = 1'b1;
	assign bitmap[2150] = 1'b0;
	assign bitmap[2151] = 1'b0;
	assign bitmap[2152] = 1'b0;
	assign bitmap[2153] = 1'b0;
	assign bitmap[2154] = 1'b1;
	assign bitmap[2155] = 1'b1;
	assign bitmap[2156] = 1'b1;
	assign bitmap[2157] = 1'b1;
	assign bitmap[2158] = 1'b0;
	assign bitmap[2159] = 1'b0;
	assign bitmap[2160] = 1'b0;
	assign bitmap[2161] = 1'b0;
	assign bitmap[2162] = 1'b0;
	assign bitmap[2163] = 1'b0;
	assign bitmap[2164] = 1'b0;
	assign bitmap[2165] = 1'b0;
	assign bitmap[2166] = 1'b0;
	assign bitmap[2167] = 1'b0;
	assign bitmap[2168] = 1'b0;
	assign bitmap[2169] = 1'b0;
	assign bitmap[2170] = 1'b0;
	assign bitmap[2171] = 1'b0;
	assign bitmap[2172] = 1'b0;
	assign bitmap[2173] = 1'b0;
	assign bitmap[2174] = 1'b0;
	assign bitmap[2175] = 1'b0;
	assign bitmap[2176] = 1'b0;
	assign bitmap[2177] = 1'b0;
	assign bitmap[2178] = 1'b0;
	assign bitmap[2179] = 1'b0;
	assign bitmap[2180] = 1'b0;
	assign bitmap[2181] = 1'b0;
	assign bitmap[2182] = 1'b0;
	assign bitmap[2183] = 1'b0;
	assign bitmap[2184] = 1'b0;
	assign bitmap[2185] = 1'b0;
	assign bitmap[2186] = 1'b0;
	assign bitmap[2187] = 1'b0;
	assign bitmap[2188] = 1'b0;
	assign bitmap[2189] = 1'b0;
	assign bitmap[2190] = 1'b0;
	assign bitmap[2191] = 1'b0;
	assign bitmap[2192] = 1'b0;
	assign bitmap[2193] = 1'b0;
	assign bitmap[2194] = 1'b1;
	assign bitmap[2195] = 1'b1;
	assign bitmap[2196] = 1'b1;
	assign bitmap[2197] = 1'b1;
	assign bitmap[2198] = 1'b0;
	assign bitmap[2199] = 1'b0;
	assign bitmap[2200] = 1'b0;
	assign bitmap[2201] = 1'b0;
	assign bitmap[2202] = 1'b0;
	assign bitmap[2203] = 1'b0;
	assign bitmap[2204] = 1'b0;
	assign bitmap[2205] = 1'b0;
	assign bitmap[2206] = 1'b0;
	assign bitmap[2207] = 1'b0;
	assign bitmap[2208] = 1'b0;
	assign bitmap[2209] = 1'b0;
	assign bitmap[2210] = 1'b1;
	assign bitmap[2211] = 1'b0;
	assign bitmap[2212] = 1'b0;
	assign bitmap[2213] = 1'b0;
	assign bitmap[2214] = 1'b0;
	assign bitmap[2215] = 1'b0;
	assign bitmap[2216] = 1'b0;
	assign bitmap[2217] = 1'b0;
	assign bitmap[2218] = 1'b0;
	assign bitmap[2219] = 1'b0;
	assign bitmap[2220] = 1'b0;
	assign bitmap[2221] = 1'b0;
	assign bitmap[2222] = 1'b0;
	assign bitmap[2223] = 1'b0;
	assign bitmap[2224] = 1'b0;
	assign bitmap[2225] = 1'b0;
	assign bitmap[2226] = 1'b1;
	assign bitmap[2227] = 1'b0;
	assign bitmap[2228] = 1'b0;
	assign bitmap[2229] = 1'b0;
	assign bitmap[2230] = 1'b0;
	assign bitmap[2231] = 1'b0;
	assign bitmap[2232] = 1'b0;
	assign bitmap[2233] = 1'b0;
	assign bitmap[2234] = 1'b0;
	assign bitmap[2235] = 1'b0;
	assign bitmap[2236] = 1'b0;
	assign bitmap[2237] = 1'b0;
	assign bitmap[2238] = 1'b0;
	assign bitmap[2239] = 1'b0;
	assign bitmap[2240] = 1'b0;
	assign bitmap[2241] = 1'b0;
	assign bitmap[2242] = 1'b1;
	assign bitmap[2243] = 1'b1;
	assign bitmap[2244] = 1'b1;
	assign bitmap[2245] = 1'b1;
	assign bitmap[2246] = 1'b0;
	assign bitmap[2247] = 1'b0;
	assign bitmap[2248] = 1'b0;
	assign bitmap[2249] = 1'b0;
	assign bitmap[2250] = 1'b0;
	assign bitmap[2251] = 1'b0;
	assign bitmap[2252] = 1'b0;
	assign bitmap[2253] = 1'b0;
	assign bitmap[2254] = 1'b0;
	assign bitmap[2255] = 1'b0;
	assign bitmap[2256] = 1'b0;
	assign bitmap[2257] = 1'b0;
	assign bitmap[2258] = 1'b1;
	assign bitmap[2259] = 1'b0;
	assign bitmap[2260] = 1'b0;
	assign bitmap[2261] = 1'b1;
	assign bitmap[2262] = 1'b0;
	assign bitmap[2263] = 1'b0;
	assign bitmap[2264] = 1'b0;
	assign bitmap[2265] = 1'b0;
	assign bitmap[2266] = 1'b0;
	assign bitmap[2267] = 1'b0;
	assign bitmap[2268] = 1'b0;
	assign bitmap[2269] = 1'b0;
	assign bitmap[2270] = 1'b0;
	assign bitmap[2271] = 1'b0;
	assign bitmap[2272] = 1'b0;
	assign bitmap[2273] = 1'b0;
	assign bitmap[2274] = 1'b1;
	assign bitmap[2275] = 1'b1;
	assign bitmap[2276] = 1'b1;
	assign bitmap[2277] = 1'b1;
	assign bitmap[2278] = 1'b0;
	assign bitmap[2279] = 1'b0;
	assign bitmap[2280] = 1'b0;
	assign bitmap[2281] = 1'b0;
	assign bitmap[2282] = 1'b0;
	assign bitmap[2283] = 1'b0;
	assign bitmap[2284] = 1'b0;
	assign bitmap[2285] = 1'b0;
	assign bitmap[2286] = 1'b0;
	assign bitmap[2287] = 1'b0;
	assign bitmap[2288] = 1'b0;
	assign bitmap[2289] = 1'b0;
	assign bitmap[2290] = 1'b0;
	assign bitmap[2291] = 1'b0;
	assign bitmap[2292] = 1'b0;
	assign bitmap[2293] = 1'b0;
	assign bitmap[2294] = 1'b0;
	assign bitmap[2295] = 1'b0;
	assign bitmap[2296] = 1'b0;
	assign bitmap[2297] = 1'b0;
	assign bitmap[2298] = 1'b0;
	assign bitmap[2299] = 1'b0;
	assign bitmap[2300] = 1'b0;
	assign bitmap[2301] = 1'b0;
	assign bitmap[2302] = 1'b0;
	assign bitmap[2303] = 1'b0;
	assign bitmap[2304] = 1'b0;
	assign bitmap[2305] = 1'b0;
	assign bitmap[2306] = 1'b0;
	assign bitmap[2307] = 1'b0;
	assign bitmap[2308] = 1'b0;
	assign bitmap[2309] = 1'b0;
	assign bitmap[2310] = 1'b0;
	assign bitmap[2311] = 1'b0;
	assign bitmap[2312] = 1'b0;
	assign bitmap[2313] = 1'b0;
	assign bitmap[2314] = 1'b0;
	assign bitmap[2315] = 1'b0;
	assign bitmap[2316] = 1'b0;
	assign bitmap[2317] = 1'b0;
	assign bitmap[2318] = 1'b0;
	assign bitmap[2319] = 1'b0;
	assign bitmap[2320] = 1'b0;
	assign bitmap[2321] = 1'b0;
	assign bitmap[2322] = 1'b1;
	assign bitmap[2323] = 1'b1;
	assign bitmap[2324] = 1'b1;
	assign bitmap[2325] = 1'b1;
	assign bitmap[2326] = 1'b0;
	assign bitmap[2327] = 1'b0;
	assign bitmap[2328] = 1'b0;
	assign bitmap[2329] = 1'b0;
	assign bitmap[2330] = 1'b0;
	assign bitmap[2331] = 1'b0;
	assign bitmap[2332] = 1'b1;
	assign bitmap[2333] = 1'b0;
	assign bitmap[2334] = 1'b0;
	assign bitmap[2335] = 1'b0;
	assign bitmap[2336] = 1'b0;
	assign bitmap[2337] = 1'b0;
	assign bitmap[2338] = 1'b1;
	assign bitmap[2339] = 1'b0;
	assign bitmap[2340] = 1'b0;
	assign bitmap[2341] = 1'b0;
	assign bitmap[2342] = 1'b0;
	assign bitmap[2343] = 1'b0;
	assign bitmap[2344] = 1'b0;
	assign bitmap[2345] = 1'b0;
	assign bitmap[2346] = 1'b0;
	assign bitmap[2347] = 1'b1;
	assign bitmap[2348] = 1'b1;
	assign bitmap[2349] = 1'b0;
	assign bitmap[2350] = 1'b0;
	assign bitmap[2351] = 1'b0;
	assign bitmap[2352] = 1'b0;
	assign bitmap[2353] = 1'b0;
	assign bitmap[2354] = 1'b1;
	assign bitmap[2355] = 1'b0;
	assign bitmap[2356] = 1'b0;
	assign bitmap[2357] = 1'b0;
	assign bitmap[2358] = 1'b0;
	assign bitmap[2359] = 1'b0;
	assign bitmap[2360] = 1'b0;
	assign bitmap[2361] = 1'b0;
	assign bitmap[2362] = 1'b1;
	assign bitmap[2363] = 1'b0;
	assign bitmap[2364] = 1'b1;
	assign bitmap[2365] = 1'b0;
	assign bitmap[2366] = 1'b0;
	assign bitmap[2367] = 1'b0;
	assign bitmap[2368] = 1'b0;
	assign bitmap[2369] = 1'b0;
	assign bitmap[2370] = 1'b1;
	assign bitmap[2371] = 1'b1;
	assign bitmap[2372] = 1'b1;
	assign bitmap[2373] = 1'b1;
	assign bitmap[2374] = 1'b0;
	assign bitmap[2375] = 1'b0;
	assign bitmap[2376] = 1'b0;
	assign bitmap[2377] = 1'b0;
	assign bitmap[2378] = 1'b0;
	assign bitmap[2379] = 1'b0;
	assign bitmap[2380] = 1'b1;
	assign bitmap[2381] = 1'b0;
	assign bitmap[2382] = 1'b0;
	assign bitmap[2383] = 1'b0;
	assign bitmap[2384] = 1'b0;
	assign bitmap[2385] = 1'b0;
	assign bitmap[2386] = 1'b0;
	assign bitmap[2387] = 1'b0;
	assign bitmap[2388] = 1'b0;
	assign bitmap[2389] = 1'b1;
	assign bitmap[2390] = 1'b0;
	assign bitmap[2391] = 1'b0;
	assign bitmap[2392] = 1'b0;
	assign bitmap[2393] = 1'b0;
	assign bitmap[2394] = 1'b0;
	assign bitmap[2395] = 1'b0;
	assign bitmap[2396] = 1'b1;
	assign bitmap[2397] = 1'b0;
	assign bitmap[2398] = 1'b0;
	assign bitmap[2399] = 1'b0;
	assign bitmap[2400] = 1'b0;
	assign bitmap[2401] = 1'b0;
	assign bitmap[2402] = 1'b1;
	assign bitmap[2403] = 1'b1;
	assign bitmap[2404] = 1'b1;
	assign bitmap[2405] = 1'b1;
	assign bitmap[2406] = 1'b0;
	assign bitmap[2407] = 1'b0;
	assign bitmap[2408] = 1'b0;
	assign bitmap[2409] = 1'b0;
	assign bitmap[2410] = 1'b1;
	assign bitmap[2411] = 1'b1;
	assign bitmap[2412] = 1'b1;
	assign bitmap[2413] = 1'b1;
	assign bitmap[2414] = 1'b0;
	assign bitmap[2415] = 1'b0;
	assign bitmap[2416] = 1'b0;
	assign bitmap[2417] = 1'b0;
	assign bitmap[2418] = 1'b0;
	assign bitmap[2419] = 1'b0;
	assign bitmap[2420] = 1'b0;
	assign bitmap[2421] = 1'b0;
	assign bitmap[2422] = 1'b0;
	assign bitmap[2423] = 1'b0;
	assign bitmap[2424] = 1'b0;
	assign bitmap[2425] = 1'b0;
	assign bitmap[2426] = 1'b0;
	assign bitmap[2427] = 1'b0;
	assign bitmap[2428] = 1'b0;
	assign bitmap[2429] = 1'b0;
	assign bitmap[2430] = 1'b0;
	assign bitmap[2431] = 1'b0;
	assign bitmap[2432] = 1'b0;
	assign bitmap[2433] = 1'b0;
	assign bitmap[2434] = 1'b0;
	assign bitmap[2435] = 1'b0;
	assign bitmap[2436] = 1'b0;
	assign bitmap[2437] = 1'b0;
	assign bitmap[2438] = 1'b0;
	assign bitmap[2439] = 1'b0;
	assign bitmap[2440] = 1'b0;
	assign bitmap[2441] = 1'b0;
	assign bitmap[2442] = 1'b0;
	assign bitmap[2443] = 1'b0;
	assign bitmap[2444] = 1'b0;
	assign bitmap[2445] = 1'b0;
	assign bitmap[2446] = 1'b0;
	assign bitmap[2447] = 1'b0;
	assign bitmap[2448] = 1'b0;
	assign bitmap[2449] = 1'b0;
	assign bitmap[2450] = 1'b0;
	assign bitmap[2451] = 1'b1;
	assign bitmap[2452] = 1'b1;
	assign bitmap[2453] = 1'b0;
	assign bitmap[2454] = 1'b0;
	assign bitmap[2455] = 1'b0;
	assign bitmap[2456] = 1'b0;
	assign bitmap[2457] = 1'b0;
	assign bitmap[2458] = 1'b0;
	assign bitmap[2459] = 1'b0;
	assign bitmap[2460] = 1'b0;
	assign bitmap[2461] = 1'b0;
	assign bitmap[2462] = 1'b0;
	assign bitmap[2463] = 1'b0;
	assign bitmap[2464] = 1'b0;
	assign bitmap[2465] = 1'b0;
	assign bitmap[2466] = 1'b1;
	assign bitmap[2467] = 1'b0;
	assign bitmap[2468] = 1'b0;
	assign bitmap[2469] = 1'b1;
	assign bitmap[2470] = 1'b0;
	assign bitmap[2471] = 1'b0;
	assign bitmap[2472] = 1'b0;
	assign bitmap[2473] = 1'b0;
	assign bitmap[2474] = 1'b0;
	assign bitmap[2475] = 1'b0;
	assign bitmap[2476] = 1'b0;
	assign bitmap[2477] = 1'b0;
	assign bitmap[2478] = 1'b0;
	assign bitmap[2479] = 1'b0;
	assign bitmap[2480] = 1'b0;
	assign bitmap[2481] = 1'b0;
	assign bitmap[2482] = 1'b0;
	assign bitmap[2483] = 1'b0;
	assign bitmap[2484] = 1'b0;
	assign bitmap[2485] = 1'b1;
	assign bitmap[2486] = 1'b0;
	assign bitmap[2487] = 1'b0;
	assign bitmap[2488] = 1'b0;
	assign bitmap[2489] = 1'b0;
	assign bitmap[2490] = 1'b0;
	assign bitmap[2491] = 1'b0;
	assign bitmap[2492] = 1'b0;
	assign bitmap[2493] = 1'b0;
	assign bitmap[2494] = 1'b0;
	assign bitmap[2495] = 1'b0;
	assign bitmap[2496] = 1'b0;
	assign bitmap[2497] = 1'b0;
	assign bitmap[2498] = 1'b0;
	assign bitmap[2499] = 1'b0;
	assign bitmap[2500] = 1'b1;
	assign bitmap[2501] = 1'b0;
	assign bitmap[2502] = 1'b0;
	assign bitmap[2503] = 1'b0;
	assign bitmap[2504] = 1'b0;
	assign bitmap[2505] = 1'b0;
	assign bitmap[2506] = 1'b0;
	assign bitmap[2507] = 1'b0;
	assign bitmap[2508] = 1'b0;
	assign bitmap[2509] = 1'b0;
	assign bitmap[2510] = 1'b0;
	assign bitmap[2511] = 1'b0;
	assign bitmap[2512] = 1'b0;
	assign bitmap[2513] = 1'b0;
	assign bitmap[2514] = 1'b0;
	assign bitmap[2515] = 1'b1;
	assign bitmap[2516] = 1'b0;
	assign bitmap[2517] = 1'b0;
	assign bitmap[2518] = 1'b0;
	assign bitmap[2519] = 1'b0;
	assign bitmap[2520] = 1'b0;
	assign bitmap[2521] = 1'b0;
	assign bitmap[2522] = 1'b0;
	assign bitmap[2523] = 1'b0;
	assign bitmap[2524] = 1'b0;
	assign bitmap[2525] = 1'b0;
	assign bitmap[2526] = 1'b0;
	assign bitmap[2527] = 1'b0;
	assign bitmap[2528] = 1'b0;
	assign bitmap[2529] = 1'b0;
	assign bitmap[2530] = 1'b1;
	assign bitmap[2531] = 1'b1;
	assign bitmap[2532] = 1'b1;
	assign bitmap[2533] = 1'b1;
	assign bitmap[2534] = 1'b0;
	assign bitmap[2535] = 1'b0;
	assign bitmap[2536] = 1'b0;
	assign bitmap[2537] = 1'b0;
	assign bitmap[2538] = 1'b0;
	assign bitmap[2539] = 1'b0;
	assign bitmap[2540] = 1'b0;
	assign bitmap[2541] = 1'b0;
	assign bitmap[2542] = 1'b0;
	assign bitmap[2543] = 1'b0;
	assign bitmap[2544] = 1'b0;
	assign bitmap[2545] = 1'b0;
	assign bitmap[2546] = 1'b0;
	assign bitmap[2547] = 1'b0;
	assign bitmap[2548] = 1'b0;
	assign bitmap[2549] = 1'b0;
	assign bitmap[2550] = 1'b0;
	assign bitmap[2551] = 1'b0;
	assign bitmap[2552] = 1'b0;
	assign bitmap[2553] = 1'b0;
	assign bitmap[2554] = 1'b0;
	assign bitmap[2555] = 1'b0;
	assign bitmap[2556] = 1'b0;
	assign bitmap[2557] = 1'b0;
	assign bitmap[2558] = 1'b0;
	assign bitmap[2559] = 1'b0;
	assign bitmap[2560] = 1'b0;
	assign bitmap[2561] = 1'b0;
	assign bitmap[2562] = 1'b0;
	assign bitmap[2563] = 1'b0;
	assign bitmap[2564] = 1'b0;
	assign bitmap[2565] = 1'b0;
	assign bitmap[2566] = 1'b0;
	assign bitmap[2567] = 1'b0;
	assign bitmap[2568] = 1'b0;
	assign bitmap[2569] = 1'b0;
	assign bitmap[2570] = 1'b0;
	assign bitmap[2571] = 1'b0;
	assign bitmap[2572] = 1'b0;
	assign bitmap[2573] = 1'b0;
	assign bitmap[2574] = 1'b0;
	assign bitmap[2575] = 1'b0;
	assign bitmap[2576] = 1'b0;
	assign bitmap[2577] = 1'b0;
	assign bitmap[2578] = 1'b0;
	assign bitmap[2579] = 1'b0;
	assign bitmap[2580] = 1'b1;
	assign bitmap[2581] = 1'b0;
	assign bitmap[2582] = 1'b0;
	assign bitmap[2583] = 1'b0;
	assign bitmap[2584] = 1'b0;
	assign bitmap[2585] = 1'b0;
	assign bitmap[2586] = 1'b1;
	assign bitmap[2587] = 1'b1;
	assign bitmap[2588] = 1'b1;
	assign bitmap[2589] = 1'b1;
	assign bitmap[2590] = 1'b0;
	assign bitmap[2591] = 1'b0;
	assign bitmap[2592] = 1'b0;
	assign bitmap[2593] = 1'b0;
	assign bitmap[2594] = 1'b0;
	assign bitmap[2595] = 1'b1;
	assign bitmap[2596] = 1'b1;
	assign bitmap[2597] = 1'b0;
	assign bitmap[2598] = 1'b0;
	assign bitmap[2599] = 1'b0;
	assign bitmap[2600] = 1'b0;
	assign bitmap[2601] = 1'b0;
	assign bitmap[2602] = 1'b1;
	assign bitmap[2603] = 1'b0;
	assign bitmap[2604] = 1'b0;
	assign bitmap[2605] = 1'b1;
	assign bitmap[2606] = 1'b0;
	assign bitmap[2607] = 1'b0;
	assign bitmap[2608] = 1'b0;
	assign bitmap[2609] = 1'b0;
	assign bitmap[2610] = 1'b1;
	assign bitmap[2611] = 1'b0;
	assign bitmap[2612] = 1'b1;
	assign bitmap[2613] = 1'b0;
	assign bitmap[2614] = 1'b0;
	assign bitmap[2615] = 1'b0;
	assign bitmap[2616] = 1'b0;
	assign bitmap[2617] = 1'b0;
	assign bitmap[2618] = 1'b1;
	assign bitmap[2619] = 1'b0;
	assign bitmap[2620] = 1'b0;
	assign bitmap[2621] = 1'b1;
	assign bitmap[2622] = 1'b0;
	assign bitmap[2623] = 1'b0;
	assign bitmap[2624] = 1'b0;
	assign bitmap[2625] = 1'b0;
	assign bitmap[2626] = 1'b0;
	assign bitmap[2627] = 1'b0;
	assign bitmap[2628] = 1'b1;
	assign bitmap[2629] = 1'b0;
	assign bitmap[2630] = 1'b0;
	assign bitmap[2631] = 1'b0;
	assign bitmap[2632] = 1'b0;
	assign bitmap[2633] = 1'b0;
	assign bitmap[2634] = 1'b1;
	assign bitmap[2635] = 1'b0;
	assign bitmap[2636] = 1'b0;
	assign bitmap[2637] = 1'b1;
	assign bitmap[2638] = 1'b0;
	assign bitmap[2639] = 1'b0;
	assign bitmap[2640] = 1'b0;
	assign bitmap[2641] = 1'b0;
	assign bitmap[2642] = 1'b0;
	assign bitmap[2643] = 1'b0;
	assign bitmap[2644] = 1'b1;
	assign bitmap[2645] = 1'b0;
	assign bitmap[2646] = 1'b0;
	assign bitmap[2647] = 1'b0;
	assign bitmap[2648] = 1'b0;
	assign bitmap[2649] = 1'b0;
	assign bitmap[2650] = 1'b1;
	assign bitmap[2651] = 1'b0;
	assign bitmap[2652] = 1'b0;
	assign bitmap[2653] = 1'b1;
	assign bitmap[2654] = 1'b0;
	assign bitmap[2655] = 1'b0;
	assign bitmap[2656] = 1'b0;
	assign bitmap[2657] = 1'b0;
	assign bitmap[2658] = 1'b1;
	assign bitmap[2659] = 1'b1;
	assign bitmap[2660] = 1'b1;
	assign bitmap[2661] = 1'b1;
	assign bitmap[2662] = 1'b0;
	assign bitmap[2663] = 1'b0;
	assign bitmap[2664] = 1'b0;
	assign bitmap[2665] = 1'b0;
	assign bitmap[2666] = 1'b1;
	assign bitmap[2667] = 1'b1;
	assign bitmap[2668] = 1'b1;
	assign bitmap[2669] = 1'b1;
	assign bitmap[2670] = 1'b0;
	assign bitmap[2671] = 1'b0;
	assign bitmap[2672] = 1'b0;
	assign bitmap[2673] = 1'b0;
	assign bitmap[2674] = 1'b0;
	assign bitmap[2675] = 1'b0;
	assign bitmap[2676] = 1'b0;
	assign bitmap[2677] = 1'b0;
	assign bitmap[2678] = 1'b0;
	assign bitmap[2679] = 1'b0;
	assign bitmap[2680] = 1'b0;
	assign bitmap[2681] = 1'b0;
	assign bitmap[2682] = 1'b0;
	assign bitmap[2683] = 1'b0;
	assign bitmap[2684] = 1'b0;
	assign bitmap[2685] = 1'b0;
	assign bitmap[2686] = 1'b0;
	assign bitmap[2687] = 1'b0;
	assign bitmap[2688] = 1'b0;
	assign bitmap[2689] = 1'b0;
	assign bitmap[2690] = 1'b0;
	assign bitmap[2691] = 1'b0;
	assign bitmap[2692] = 1'b0;
	assign bitmap[2693] = 1'b0;
	assign bitmap[2694] = 1'b0;
	assign bitmap[2695] = 1'b0;
	assign bitmap[2696] = 1'b0;
	assign bitmap[2697] = 1'b0;
	assign bitmap[2698] = 1'b0;
	assign bitmap[2699] = 1'b0;
	assign bitmap[2700] = 1'b0;
	assign bitmap[2701] = 1'b0;
	assign bitmap[2702] = 1'b0;
	assign bitmap[2703] = 1'b0;
	assign bitmap[2704] = 1'b0;
	assign bitmap[2705] = 1'b0;
	assign bitmap[2706] = 1'b0;
	assign bitmap[2707] = 1'b1;
	assign bitmap[2708] = 1'b1;
	assign bitmap[2709] = 1'b0;
	assign bitmap[2710] = 1'b0;
	assign bitmap[2711] = 1'b0;
	assign bitmap[2712] = 1'b0;
	assign bitmap[2713] = 1'b0;
	assign bitmap[2714] = 1'b0;
	assign bitmap[2715] = 1'b0;
	assign bitmap[2716] = 1'b1;
	assign bitmap[2717] = 1'b1;
	assign bitmap[2718] = 1'b0;
	assign bitmap[2719] = 1'b0;
	assign bitmap[2720] = 1'b0;
	assign bitmap[2721] = 1'b0;
	assign bitmap[2722] = 1'b1;
	assign bitmap[2723] = 1'b0;
	assign bitmap[2724] = 1'b0;
	assign bitmap[2725] = 1'b1;
	assign bitmap[2726] = 1'b0;
	assign bitmap[2727] = 1'b0;
	assign bitmap[2728] = 1'b0;
	assign bitmap[2729] = 1'b0;
	assign bitmap[2730] = 1'b0;
	assign bitmap[2731] = 1'b1;
	assign bitmap[2732] = 1'b0;
	assign bitmap[2733] = 1'b1;
	assign bitmap[2734] = 1'b0;
	assign bitmap[2735] = 1'b0;
	assign bitmap[2736] = 1'b0;
	assign bitmap[2737] = 1'b0;
	assign bitmap[2738] = 1'b0;
	assign bitmap[2739] = 1'b0;
	assign bitmap[2740] = 1'b0;
	assign bitmap[2741] = 1'b1;
	assign bitmap[2742] = 1'b0;
	assign bitmap[2743] = 1'b0;
	assign bitmap[2744] = 1'b0;
	assign bitmap[2745] = 1'b0;
	assign bitmap[2746] = 1'b1;
	assign bitmap[2747] = 1'b0;
	assign bitmap[2748] = 1'b0;
	assign bitmap[2749] = 1'b1;
	assign bitmap[2750] = 1'b0;
	assign bitmap[2751] = 1'b0;
	assign bitmap[2752] = 1'b0;
	assign bitmap[2753] = 1'b0;
	assign bitmap[2754] = 1'b0;
	assign bitmap[2755] = 1'b0;
	assign bitmap[2756] = 1'b1;
	assign bitmap[2757] = 1'b0;
	assign bitmap[2758] = 1'b0;
	assign bitmap[2759] = 1'b0;
	assign bitmap[2760] = 1'b0;
	assign bitmap[2761] = 1'b0;
	assign bitmap[2762] = 1'b1;
	assign bitmap[2763] = 1'b1;
	assign bitmap[2764] = 1'b1;
	assign bitmap[2765] = 1'b1;
	assign bitmap[2766] = 1'b1;
	assign bitmap[2767] = 1'b0;
	assign bitmap[2768] = 1'b0;
	assign bitmap[2769] = 1'b0;
	assign bitmap[2770] = 1'b0;
	assign bitmap[2771] = 1'b1;
	assign bitmap[2772] = 1'b0;
	assign bitmap[2773] = 1'b0;
	assign bitmap[2774] = 1'b0;
	assign bitmap[2775] = 1'b0;
	assign bitmap[2776] = 1'b0;
	assign bitmap[2777] = 1'b0;
	assign bitmap[2778] = 1'b0;
	assign bitmap[2779] = 1'b0;
	assign bitmap[2780] = 1'b0;
	assign bitmap[2781] = 1'b1;
	assign bitmap[2782] = 1'b0;
	assign bitmap[2783] = 1'b0;
	assign bitmap[2784] = 1'b0;
	assign bitmap[2785] = 1'b0;
	assign bitmap[2786] = 1'b1;
	assign bitmap[2787] = 1'b1;
	assign bitmap[2788] = 1'b1;
	assign bitmap[2789] = 1'b1;
	assign bitmap[2790] = 1'b0;
	assign bitmap[2791] = 1'b0;
	assign bitmap[2792] = 1'b0;
	assign bitmap[2793] = 1'b0;
	assign bitmap[2794] = 1'b0;
	assign bitmap[2795] = 1'b0;
	assign bitmap[2796] = 1'b0;
	assign bitmap[2797] = 1'b1;
	assign bitmap[2798] = 1'b0;
	assign bitmap[2799] = 1'b0;
	assign bitmap[2800] = 1'b0;
	assign bitmap[2801] = 1'b0;
	assign bitmap[2802] = 1'b0;
	assign bitmap[2803] = 1'b0;
	assign bitmap[2804] = 1'b0;
	assign bitmap[2805] = 1'b0;
	assign bitmap[2806] = 1'b0;
	assign bitmap[2807] = 1'b0;
	assign bitmap[2808] = 1'b0;
	assign bitmap[2809] = 1'b0;
	assign bitmap[2810] = 1'b0;
	assign bitmap[2811] = 1'b0;
	assign bitmap[2812] = 1'b0;
	assign bitmap[2813] = 1'b0;
	assign bitmap[2814] = 1'b0;
	assign bitmap[2815] = 1'b0;
	assign bitmap[2816] = 1'b0;
	assign bitmap[2817] = 1'b0;
	assign bitmap[2818] = 1'b0;
	assign bitmap[2819] = 1'b0;
	assign bitmap[2820] = 1'b0;
	assign bitmap[2821] = 1'b0;
	assign bitmap[2822] = 1'b0;
	assign bitmap[2823] = 1'b0;
	assign bitmap[2824] = 1'b0;
	assign bitmap[2825] = 1'b0;
	assign bitmap[2826] = 1'b0;
	assign bitmap[2827] = 1'b0;
	assign bitmap[2828] = 1'b0;
	assign bitmap[2829] = 1'b0;
	assign bitmap[2830] = 1'b0;
	assign bitmap[2831] = 1'b0;
	assign bitmap[2832] = 1'b0;
	assign bitmap[2833] = 1'b0;
	assign bitmap[2834] = 1'b0;
	assign bitmap[2835] = 1'b1;
	assign bitmap[2836] = 1'b1;
	assign bitmap[2837] = 1'b0;
	assign bitmap[2838] = 1'b0;
	assign bitmap[2839] = 1'b0;
	assign bitmap[2840] = 1'b0;
	assign bitmap[2841] = 1'b0;
	assign bitmap[2842] = 1'b1;
	assign bitmap[2843] = 1'b1;
	assign bitmap[2844] = 1'b1;
	assign bitmap[2845] = 1'b1;
	assign bitmap[2846] = 1'b0;
	assign bitmap[2847] = 1'b0;
	assign bitmap[2848] = 1'b0;
	assign bitmap[2849] = 1'b0;
	assign bitmap[2850] = 1'b1;
	assign bitmap[2851] = 1'b0;
	assign bitmap[2852] = 1'b0;
	assign bitmap[2853] = 1'b1;
	assign bitmap[2854] = 1'b0;
	assign bitmap[2855] = 1'b0;
	assign bitmap[2856] = 1'b0;
	assign bitmap[2857] = 1'b0;
	assign bitmap[2858] = 1'b1;
	assign bitmap[2859] = 1'b0;
	assign bitmap[2860] = 1'b0;
	assign bitmap[2861] = 1'b1;
	assign bitmap[2862] = 1'b0;
	assign bitmap[2863] = 1'b0;
	assign bitmap[2864] = 1'b0;
	assign bitmap[2865] = 1'b0;
	assign bitmap[2866] = 1'b0;
	assign bitmap[2867] = 1'b0;
	assign bitmap[2868] = 1'b0;
	assign bitmap[2869] = 1'b1;
	assign bitmap[2870] = 1'b0;
	assign bitmap[2871] = 1'b0;
	assign bitmap[2872] = 1'b0;
	assign bitmap[2873] = 1'b0;
	assign bitmap[2874] = 1'b1;
	assign bitmap[2875] = 1'b0;
	assign bitmap[2876] = 1'b0;
	assign bitmap[2877] = 1'b1;
	assign bitmap[2878] = 1'b0;
	assign bitmap[2879] = 1'b0;
	assign bitmap[2880] = 1'b0;
	assign bitmap[2881] = 1'b0;
	assign bitmap[2882] = 1'b0;
	assign bitmap[2883] = 1'b0;
	assign bitmap[2884] = 1'b1;
	assign bitmap[2885] = 1'b0;
	assign bitmap[2886] = 1'b0;
	assign bitmap[2887] = 1'b0;
	assign bitmap[2888] = 1'b0;
	assign bitmap[2889] = 1'b0;
	assign bitmap[2890] = 1'b1;
	assign bitmap[2891] = 1'b0;
	assign bitmap[2892] = 1'b0;
	assign bitmap[2893] = 1'b1;
	assign bitmap[2894] = 1'b0;
	assign bitmap[2895] = 1'b0;
	assign bitmap[2896] = 1'b0;
	assign bitmap[2897] = 1'b0;
	assign bitmap[2898] = 1'b0;
	assign bitmap[2899] = 1'b1;
	assign bitmap[2900] = 1'b0;
	assign bitmap[2901] = 1'b0;
	assign bitmap[2902] = 1'b0;
	assign bitmap[2903] = 1'b0;
	assign bitmap[2904] = 1'b0;
	assign bitmap[2905] = 1'b0;
	assign bitmap[2906] = 1'b1;
	assign bitmap[2907] = 1'b0;
	assign bitmap[2908] = 1'b0;
	assign bitmap[2909] = 1'b1;
	assign bitmap[2910] = 1'b0;
	assign bitmap[2911] = 1'b0;
	assign bitmap[2912] = 1'b0;
	assign bitmap[2913] = 1'b0;
	assign bitmap[2914] = 1'b1;
	assign bitmap[2915] = 1'b1;
	assign bitmap[2916] = 1'b1;
	assign bitmap[2917] = 1'b1;
	assign bitmap[2918] = 1'b0;
	assign bitmap[2919] = 1'b0;
	assign bitmap[2920] = 1'b0;
	assign bitmap[2921] = 1'b0;
	assign bitmap[2922] = 1'b1;
	assign bitmap[2923] = 1'b1;
	assign bitmap[2924] = 1'b1;
	assign bitmap[2925] = 1'b1;
	assign bitmap[2926] = 1'b0;
	assign bitmap[2927] = 1'b0;
	assign bitmap[2928] = 1'b0;
	assign bitmap[2929] = 1'b0;
	assign bitmap[2930] = 1'b0;
	assign bitmap[2931] = 1'b0;
	assign bitmap[2932] = 1'b0;
	assign bitmap[2933] = 1'b0;
	assign bitmap[2934] = 1'b0;
	assign bitmap[2935] = 1'b0;
	assign bitmap[2936] = 1'b0;
	assign bitmap[2937] = 1'b0;
	assign bitmap[2938] = 1'b0;
	assign bitmap[2939] = 1'b0;
	assign bitmap[2940] = 1'b0;
	assign bitmap[2941] = 1'b0;
	assign bitmap[2942] = 1'b0;
	assign bitmap[2943] = 1'b0;
	assign bitmap[2944] = 1'b0;
	assign bitmap[2945] = 1'b0;
	assign bitmap[2946] = 1'b0;
	assign bitmap[2947] = 1'b0;
	assign bitmap[2948] = 1'b0;
	assign bitmap[2949] = 1'b0;
	assign bitmap[2950] = 1'b0;
	assign bitmap[2951] = 1'b0;
	assign bitmap[2952] = 1'b0;
	assign bitmap[2953] = 1'b0;
	assign bitmap[2954] = 1'b0;
	assign bitmap[2955] = 1'b0;
	assign bitmap[2956] = 1'b0;
	assign bitmap[2957] = 1'b0;
	assign bitmap[2958] = 1'b0;
	assign bitmap[2959] = 1'b0;
	assign bitmap[2960] = 1'b0;
	assign bitmap[2961] = 1'b0;
	assign bitmap[2962] = 1'b0;
	assign bitmap[2963] = 1'b0;
	assign bitmap[2964] = 1'b1;
	assign bitmap[2965] = 1'b1;
	assign bitmap[2966] = 1'b0;
	assign bitmap[2967] = 1'b0;
	assign bitmap[2968] = 1'b0;
	assign bitmap[2969] = 1'b0;
	assign bitmap[2970] = 1'b1;
	assign bitmap[2971] = 1'b1;
	assign bitmap[2972] = 1'b1;
	assign bitmap[2973] = 1'b1;
	assign bitmap[2974] = 1'b0;
	assign bitmap[2975] = 1'b0;
	assign bitmap[2976] = 1'b0;
	assign bitmap[2977] = 1'b0;
	assign bitmap[2978] = 1'b0;
	assign bitmap[2979] = 1'b1;
	assign bitmap[2980] = 1'b0;
	assign bitmap[2981] = 1'b1;
	assign bitmap[2982] = 1'b0;
	assign bitmap[2983] = 1'b0;
	assign bitmap[2984] = 1'b0;
	assign bitmap[2985] = 1'b0;
	assign bitmap[2986] = 1'b1;
	assign bitmap[2987] = 1'b0;
	assign bitmap[2988] = 1'b0;
	assign bitmap[2989] = 1'b1;
	assign bitmap[2990] = 1'b0;
	assign bitmap[2991] = 1'b0;
	assign bitmap[2992] = 1'b0;
	assign bitmap[2993] = 1'b0;
	assign bitmap[2994] = 1'b1;
	assign bitmap[2995] = 1'b0;
	assign bitmap[2996] = 1'b0;
	assign bitmap[2997] = 1'b1;
	assign bitmap[2998] = 1'b0;
	assign bitmap[2999] = 1'b0;
	assign bitmap[3000] = 1'b0;
	assign bitmap[3001] = 1'b0;
	assign bitmap[3002] = 1'b1;
	assign bitmap[3003] = 1'b0;
	assign bitmap[3004] = 1'b0;
	assign bitmap[3005] = 1'b1;
	assign bitmap[3006] = 1'b0;
	assign bitmap[3007] = 1'b0;
	assign bitmap[3008] = 1'b0;
	assign bitmap[3009] = 1'b0;
	assign bitmap[3010] = 1'b1;
	assign bitmap[3011] = 1'b1;
	assign bitmap[3012] = 1'b1;
	assign bitmap[3013] = 1'b1;
	assign bitmap[3014] = 1'b1;
	assign bitmap[3015] = 1'b0;
	assign bitmap[3016] = 1'b0;
	assign bitmap[3017] = 1'b0;
	assign bitmap[3018] = 1'b1;
	assign bitmap[3019] = 1'b1;
	assign bitmap[3020] = 1'b1;
	assign bitmap[3021] = 1'b1;
	assign bitmap[3022] = 1'b0;
	assign bitmap[3023] = 1'b0;
	assign bitmap[3024] = 1'b0;
	assign bitmap[3025] = 1'b0;
	assign bitmap[3026] = 1'b0;
	assign bitmap[3027] = 1'b0;
	assign bitmap[3028] = 1'b0;
	assign bitmap[3029] = 1'b1;
	assign bitmap[3030] = 1'b0;
	assign bitmap[3031] = 1'b0;
	assign bitmap[3032] = 1'b0;
	assign bitmap[3033] = 1'b0;
	assign bitmap[3034] = 1'b1;
	assign bitmap[3035] = 1'b0;
	assign bitmap[3036] = 1'b0;
	assign bitmap[3037] = 1'b1;
	assign bitmap[3038] = 1'b0;
	assign bitmap[3039] = 1'b0;
	assign bitmap[3040] = 1'b0;
	assign bitmap[3041] = 1'b0;
	assign bitmap[3042] = 1'b0;
	assign bitmap[3043] = 1'b0;
	assign bitmap[3044] = 1'b0;
	assign bitmap[3045] = 1'b1;
	assign bitmap[3046] = 1'b0;
	assign bitmap[3047] = 1'b0;
	assign bitmap[3048] = 1'b0;
	assign bitmap[3049] = 1'b0;
	assign bitmap[3050] = 1'b1;
	assign bitmap[3051] = 1'b1;
	assign bitmap[3052] = 1'b1;
	assign bitmap[3053] = 1'b1;
	assign bitmap[3054] = 1'b0;
	assign bitmap[3055] = 1'b0;
	assign bitmap[3056] = 1'b0;
	assign bitmap[3057] = 1'b0;
	assign bitmap[3058] = 1'b0;
	assign bitmap[3059] = 1'b0;
	assign bitmap[3060] = 1'b0;
	assign bitmap[3061] = 1'b0;
	assign bitmap[3062] = 1'b0;
	assign bitmap[3063] = 1'b0;
	assign bitmap[3064] = 1'b0;
	assign bitmap[3065] = 1'b0;
	assign bitmap[3066] = 1'b0;
	assign bitmap[3067] = 1'b0;
	assign bitmap[3068] = 1'b0;
	assign bitmap[3069] = 1'b0;
	assign bitmap[3070] = 1'b0;
	assign bitmap[3071] = 1'b0;

	assign palette[0]  = 12'b1111_1111_1111;
	assign palette[1]  = 12'b0000_0000_0000;
	assign palette[2]  = 12'b1111_0000_0000;
	assign palette[3]  = 12'b0000_0000_0000;
	assign palette[4]  = 12'b1111_1000_0000;
	assign palette[5]  = 12'b0000_0000_0000;
	assign palette[6]  = 12'b1111_1111_0000;
	assign palette[7]  = 12'b0000_0000_0000;
	assign palette[8]  = 12'b1000_1111_0000;
	assign palette[9]  = 12'b0000_0000_0000;
	assign palette[10] = 12'b0000_1111_0000;
	assign palette[11] = 12'b0000_0000_0000;
	assign palette[12] = 12'b0000_1111_1000;
	assign palette[13] = 12'b0000_0000_0000;
	assign palette[14] = 12'b0000_1111_1111;
	assign palette[15] = 12'b0000_0000_0000;
	assign palette[16] = 12'b0000_1000_1111;
	assign palette[17] = 12'b0000_0000_0000;
	assign palette[18] = 12'b0000_0000_1111;
	assign palette[19] = 12'b0000_0000_0000;
	assign palette[20] = 12'b1000_0000_1111;
	assign palette[21] = 12'b0000_0000_0000;
	assign palette[22] = 12'b1111_0000_1111;
	assign palette[23] = 12'b0000_0000_0000;

endmodule
