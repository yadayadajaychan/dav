module miniALU (
    // TODO: define your input and output ports

    );

    // The following block contains the logic of your combinational circuit
    always_comb begin
        // TODO: write the logic for your miniALU here

    end
endmodule