module miniALU_top (
	// TODO: define your input and output ports
	input [9:0] in,
	output [9:0] out
);
    assign out = in;
endmodule
